library ieee;
use ieee.std_logic_1164.all;

--
--package common is
--
--	type pic_array is array(0 downto 4799) of std_logic;
--	
--end common;
--
--package body common is 
--end common;
--
entity Display_Frame is
--	--type pic_array is array(0 downto 4799) of std_logic;
--	Port (cont_pic : out pic_array);
--	
end entity;
--
--
architecture Display_Arc of Display_Frame is 
--
--	
--	signal Constant_pic : pic_array;
--	
	begin
--	
--	
end architecture;