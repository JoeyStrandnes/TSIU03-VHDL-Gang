library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pixel_reg is
  Port ( clk, rstn     : in std_logic;
         up_lo_byte    : in std_logic; -- '0' <=> read lo byte.
         pixcode       : out unsigned(7 downto 0);
         -- RAM signals
         --Constant_pic : in std_logic;
			higher_byte, lower_byte : in unsigned(7 downto 0));
			
end entity;

architecture rtl of pixel_reg is


type pic_array is array(0 to 4799) of std_logic;
signal Constant_pic : pic_array;
signal row, col :  unsigned(6 downto 0);
signal index : integer;

begin
	Constant_pic <= ('0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1');
	process(clk)
	begin
		if (rising_edge(clk)) then
			
			for vert in 0 to 59 loop
			
				for upscale_y in 0 to 7 loop
			
					for hort in 0 to 79 loop
			
						for upscale_x in 0 to 7 loop
								
							pixcode <= "10001100";
							--index <= to_integer(row*60 + col);
							--pixcode <= "1000000" & Constant_pic(index); --row*60 + col
							--pixcode <= Constant_pic(to_unsigned(60, (7 downto 0)));
							
						end loop;
						col <= col+1;
					end loop;
					col <= "0000000";
				end loop;
				row <= row+1;
			end loop;
			row <= "0000000";
			
			
			
--			if (up_lo_byte = '1') then
--				pixcode <= higher_byte;
--			else
--				pixcode <= lower_byte;				
--			end if;
		end if;
	end process;

end architecture;
