library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity wavefile is
  port(clk  : in std_logic;
       addr : in unsigned(13-1 downto 0); -- range 0..6470-1
       data : out signed(16-1 downto 0)); -- latency=2 clock cycles
end entity;

architecture rtl of wavefile is
  constant Nrows : integer := 6470; -- total size
  constant NBlockAbits : integer := 10; -- Each block has 2^NBlockAbits
  constant NBlocks : integer := (Nrows-1)/2**NBlockAbits+1; -- = 7
  -- Strategy:
  -- Implement NBlocks number of M9k memories (2^NBlockAbits x 9 bits).
  -- Declare a small array of length NBlocks, where each element is the output from an M9k.
  -- Put a (registered) multiplexer on the output.
  subtype word_t is signed(9-1 downto 0);
  type m9k_t is array(0 to 2**NBlockAbits-1) of word_t;
  type rom_out_vec_t is array(0 to NBlocks-1) of word_t;
  signal data_vec : rom_out_vec_t; -- assigned from NBlocks different ROMs.
  signal rom0,rom1,rom2,rom3,rom4,rom5,rom6 : m9k_t;
  signal addr_upper : unsigned(addr'left-NBlockAbits downto 0);
begin
  process(clk) begin
    if rising_edge(clk) then
      -- Generate the NBlocks M9k memories (pipelined output):
      data_vec(0) <= rom0(to_integer(addr(NBlockAbits-1 downto 0)));
      data_vec(1) <= rom1(to_integer(addr(NBlockAbits-1 downto 0)));
      data_vec(2) <= rom2(to_integer(addr(NBlockAbits-1 downto 0)));
      data_vec(3) <= rom3(to_integer(addr(NBlockAbits-1 downto 0)));
      data_vec(4) <= rom4(to_integer(addr(NBlockAbits-1 downto 0)));
      data_vec(5) <= rom5(to_integer(addr(NBlockAbits-1 downto 0)));
      data_vec(6) <= rom6(to_integer(addr(NBlockAbits-1 downto 0)));
      -- Also pipeline the upper part of the address:
      addr_upper <= addr(addr'left downto NBlockAbits);
      
      -- Use the upper address to multiplex the right output:
      data <= data_vec(to_integer(addr_upper));
    end if;
  end process;
  
  -- Last thing to do: Define the content of rom<0..6>:
  rom0 <= (
0=>"0101101000010000",
1=>"0110110010001101",
2=>"1110100010111010",
3=>"1011100100111000",
4=>"1101110100010110",
5=>"0001110100010110",
6=>"0001110100101100",
7=>"1110100010011111",
8=>"1101101110101111",
9=>"0000000011110011",
10=>"0001001100001010",
11=>"0000111000001110",
12=>"1100110010101101",
13=>"1100010010010000",
14=>"0100010011001111",
15=>"0111100110000101",
16=>"0000100010001101",
17=>"1011100101000001",
18=>"1101000001010100",
19=>"0000111110101110",
20=>"0010010011000010",
21=>"1111010000110110",
22=>"1101100010001101",
23=>"1111100011110111",
24=>"0001000001011110",
25=>"0001001110000001",
26=>"1101110111100110",
27=>"1011011100001000",
28=>"0010001001011001",
29=>"0111111111111111",
30=>"0010100001111001",
31=>"1100000011111000",
32=>"1100010100001011",
33=>"0000000100100101",
34=>"0010100000011111",
35=>"0000001101011101",
36=>"1101011111100000",
37=>"1110111110111111",
38=>"0000110011011001",
39=>"0001010111011010",
40=>"1111000000000001",
41=>"1011010100110000",
42=>"1111111100101001",
43=>"0111101000011110",
44=>"0100011010111001",
45=>"1101000001110001",
46=>"1011101111011101",
47=>"1111000111001011",
48=>"0010010000111001",
49=>"0001000101100101",
50=>"1101110001010010",
51=>"1110011001000101",
52=>"0000011111010100",
53=>"0001010111100111",
54=>"1111111011000010",
55=>"1011110001000100",
56=>"1101111101101000",
57=>"0110011110110011",
58=>"0110001001110110",
59=>"1110010111100111",
60=>"1011011111010100",
61=>"1110001010011001",
62=>"0001110010101000",
63=>"0001110000000110",
64=>"1110010100000010",
65=>"1101111011011100",
66=>"0000000111110011",
67=>"0001010001011101",
68=>"0000101010100100",
69=>"1100101000000100",
70=>"1100100000000111",
71=>"0100110001110110",
72=>"0111011010010111",
73=>"0000001001011010",
74=>"1011011101000001",
75=>"1101001111011111",
76=>"0001001011001010",
77=>"0010010000010110",
78=>"1111000011110010",
79=>"1101100101100110",
80=>"1111101001101100",
81=>"0001001000001000",
82=>"0001001000100110",
83=>"1101101001111100",
84=>"1011100011000000",
85=>"0010101100101010",
86=>"0111111011101101",
87=>"0010000100100101",
88=>"1011111011100011",
89=>"1100011110010110",
90=>"0000001110111110",
91=>"0010100000101000",
92=>"1111111100111011",
93=>"1101011110111001",
94=>"1111000100100100",
95=>"0000111010101100",
96=>"0001010100110110",
97=>"1110110010010011",
98=>"1011010011010000",
99=>"0000011011011111",
100=>"0111101110101001",
101=>"0100000010110111",
102=>"1100110000011111",
103=>"1011110110101011",
104=>"1111010100111001",
105=>"0010011001001100",
106=>"0000110101110010",
107=>"1101110000000011",
108=>"1110011001010100",
109=>"0000100100000000",
110=>"0001011000010010",
111=>"1111111001010101",
112=>"1011101011011010",
113=>"1110000110000101",
114=>"0110100010000111",
115=>"0110000110111000",
116=>"1110010110100110",
117=>"1011011100100101",
118=>"1110001111100101",
119=>"0001110100110111",
120=>"0001101111100000",
121=>"1110001111110001",
122=>"1101111011100100",
123=>"0000001000110010",
124=>"0001010000010111",
125=>"0000101010001001",
126=>"1100011111101111",
127=>"1100100011000001",
128=>"0100110110001101",
129=>"0111010101000111",
130=>"0000000011010010",
131=>"1011011110110011",
132=>"1101010010111011",
133=>"0001001001110111",
134=>"0010001111100011",
135=>"1111000010111111",
136=>"1101100100110011",
137=>"1111101100110111",
138=>"0001000110101100",
139=>"0001000101110111",
140=>"1101100101101011",
141=>"1011101000001101",
142=>"0010110000111000",
143=>"0111111010100010",
144=>"0001111101001111",
145=>"1011111000100111",
146=>"1100100000010101",
147=>"0000010101001011",
148=>"0010011110101010",
149=>"1111111101011111",
150=>"1101011110001010",
151=>"1111000111111010",
152=>"0000111010100101",
153=>"0001010100011111",
154=>"1110101101000010",
155=>"1011010100010001",
156=>"0000100010001110",
157=>"0111110010011110",
158=>"0011111011010011",
159=>"1100101110111010",
160=>"1011111001101001",
161=>"1111011001011110",
162=>"0010011001010010",
163=>"0000110011110110",
164=>"1101101000110101",
165=>"1110100001101000",
166=>"0000100011101100",
167=>"0001011000101101",
168=>"1111101101110101",
169=>"1011100101011011",
170=>"1110100000111001",
171=>"0110110111001011",
172=>"0101110000010111",
173=>"1101111110011100",
174=>"1011011111001010",
175=>"1110011011011100",
176=>"0001111110011111",
177=>"0001100100101001",
178=>"1110001001000000",
179=>"1110000000011100",
180=>"0000010000010000",
181=>"0001001111111101",
182=>"0000100001000001",
183=>"1100010011001111",
184=>"1100110110100010",
185=>"0101010010110111",
186=>"0111001000010000",
187=>"1111101000000010",
188=>"1011011100000010",
189=>"1101100001100001",
190=>"0001010011100111",
191=>"0010001011100111",
192=>"1110111000000011",
193=>"1101101010100000",
194=>"1111110010110100",
195=>"0001001000110000",
196=>"0001000010001100",
197=>"1101010111011001",
198=>"1011110001110101",
199=>"0011010001000110",
200=>"0111110110010010",
201=>"0001100010001110",
202=>"1011110001101111",
203=>"1100101011000100",
204=>"0000100001110101",
205=>"0010011011101000",
206=>"1111101110101001",
207=>"1101011110010011",
208=>"1111001111100001",
209=>"0000111101110011",
210=>"0001010100000001",
211=>"1110011011001010",
212=>"1011010101000011",
213=>"0000110001110101",
214=>"0111110001100011",
215=>"0011110101001101",
216=>"1100100111111011",
217=>"1011111110000000",
218=>"1111011010010011",
219=>"0010010111010101",
220=>"0000101110101100",
221=>"1101101011000010",
222=>"1110100101110001",
223=>"0000101000010110",
224=>"0001010111111100",
225=>"1111101011010011",
226=>"1011100100110111",
227=>"1110101000110100",
228=>"0110111100000111",
229=>"0101101011101010",
230=>"1101111000110000",
231=>"1011011111011110",
232=>"1110011110100010",
233=>"0010000011011101",
234=>"0001100000110000",
235=>"1110000111000110",
236=>"1110000011011010",
237=>"0000010010100000",
238=>"0001010100111010",
239=>"0000011110100101",
240=>"1100001111100110",
241=>"1100111100000110",
242=>"0101011010010100",
243=>"0111000010011000",
244=>"1111100000100100",
245=>"1011011110010010",
246=>"1101100000111100",
247=>"0001011000001100",
248=>"0010001010001100",
249=>"1110110010110101",
250=>"1101101001001011",
251=>"1111110100010010",
252=>"0001001100010101",
253=>"0000111110110100",
254=>"1101010100000100",
255=>"1011110011000110",
256=>"0011010111011101",
257=>"0111110101010101",
258=>"0001011001011010",
259=>"1011101110010110",
260=>"1100101100011011",
261=>"0000100110001110",
262=>"0010011100110110",
263=>"1111101010000101",
264=>"1101011110100001",
265=>"1111010000010111",
266=>"0000111100110001",
267=>"0001010100101001",
268=>"1110011100000011",
269=>"1011010100111011",
270=>"0001001101100110",
271=>"0111111000101111",
272=>"0011011010011010",
273=>"1100011100011011",
274=>"1100000001100100",
275=>"1111101001010010",
276=>"0010011011010000",
277=>"0000100001101111",
278=>"1101100110001000",
279=>"1110101110111111",
280=>"0000101011101000",
281=>"0001011000111000",
282=>"1111011100011000",
283=>"1011011010000100",
284=>"1111000010111000",
285=>"0111001100001010",
286=>"0101010011011100",
287=>"1101100100001000",
288=>"1011100110000101",
289=>"1110101011100111",
290=>"0010001000111101",
291=>"0001011100010011",
292=>"1101111110100000",
293=>"1110001011000110",
294=>"0000010110011001",
295=>"0001010101010010",
296=>"0000010010111000",
297=>"1100000101111100",
298=>"1101001111000000",
299=>"0101110100000111",
300=>"0110110000010111",
301=>"1111000110110010",
302=>"1011011011100011",
303=>"1101101110111010",
304=>"0001100001011100",
305=>"0010000010110101",
306=>"1110101010010010",
307=>"1101101101111001",
308=>"1111111010010011",
309=>"0001001100000001",
310=>"0000111000011100",
311=>"1101000010111110",
312=>"1011111111101011",
313=>"0011110101001001",
314=>"0111101111001111",
315=>"0000111011001111",
316=>"1011101001110011",
317=>"1100111001100011",
318=>"0000110000010101",
319=>"0010010110001010",
320=>"1111100010111011",
321=>"1101011110101111",
322=>"1111010001001100",
323=>"0000111100000111",
324=>"0001010010011111",
325=>"1110010110011011",
326=>"1011010101001111",
327=>"0001010011101110",
328=>"0111111010111100",
329=>"0011010100000110",
330=>"1100010111110010",
331=>"1100000011011101",
332=>"1111101110000111",
333=>"0010011010110000",
334=>"0000100000110110",
335=>"1101100100000001",
336=>"1110101111001000",
337=>"0000101100101111",
338=>"0001010101101010",
339=>"1111011011000111",
340=>"1011011000101101",
341=>"1111001011111011",
342=>"0111001111001111",
343=>"0101001101100010",
344=>"1101011111010000",
345=>"1011101000001010",
346=>"1110101111011110",
347=>"0010000111011011",
348=>"0001011000011001",
349=>"1101111110001101",
350=>"1110001101100000",
351=>"0000010111101010",
352=>"0001010101001111",
353=>"0000010001110111",
354=>"1100000011000000",
355=>"1101010111100011",
356=>"0101110111001110",
357=>"0110101100111110",
358=>"1111000011001101",
359=>"1011011100100111",
360=>"1101110010110111",
361=>"0001100101001000",
362=>"0001111111001111",
363=>"1110100110110011",
364=>"1101101110110100",
365=>"1111111100111000",
366=>"0001001111010101",
367=>"0000110110111111",
368=>"1100111110000011",
369=>"1100000010000000",
370=>"0011111110001100",
371=>"0111101010111101",
372=>"0000111011101101",
373=>"1011100101010110",
374=>"1100111101011110",
375=>"0000110011011000",
376=>"0010010111101011",
377=>"1111011001110100",
378=>"1101011111000110",
379=>"1111011100111010",
380=>"0000111110100100",
381=>"0001010000101011",
382=>"1110000100011101",
383=>"1011010111100000",
384=>"0001110010011000",
385=>"0111111100000110",
386=>"0010110111111100",
387=>"1100001101001111",
388=>"1100001100110111",
389=>"1111111001111100",
390=>"0010011100001011",
391=>"0000010101101100",
392=>"1101100000111100",
393=>"1110111001000001",
394=>"0000110001101110",
395=>"0001010111011100",
396=>"1111001001111101",
397=>"1011010111111111",
398=>"1111100111101001",
399=>"0111011011110110",
400=>"0100110000111000",
401=>"1101001110001100",
402=>"1011101011111101",
403=>"1110111101011011",
404=>"0010001111000111",
405=>"0001001101111011",
406=>"1101110110011100",
407=>"1110010010101001",
408=>"0000011110101010",
409=>"0001010111011000",
410=>"0000000100000001",
411=>"1011111001001011",
412=>"1101101011111101",
413=>"0110001110111110",
414=>"0110011001101110",
415=>"1110101010011111",
416=>"1011011101101100",
417=>"1110000000011010",
418=>"0001110000000010",
419=>"0001111000110000",
420=>"1110011001110110",
421=>"1101110011111111",
422=>"0000000000010010",
423=>"0001001110111011",
424=>"0000110000111010",
425=>"1100110001111100",
426=>"1100001011010111",
427=>"0100000110011001",
428=>"0111101001100010",
429=>"0000110001001101",
430=>"1011100101110011",
431=>"1100111101000111",
432=>"0000110111011011",
433=>"0010010110011011",
434=>"1111010101100000",
435=>"1101100010011101",
436=>"1111011110110111",
437=>"0001000001001101",
438=>"0001001110101011",
439=>"1110000000101100",
440=>"1011011000000010",
441=>"0001111010111100",
442=>"0111111110101011",
443=>"0010110000111101",
444=>"1100001000001001",
445=>"1100010000100101",
446=>"1111111101000111",
447=>"0010100001000000",
448=>"0000010010111111",
449=>"1101100001010011",
450=>"1110111010000111",
451=>"0000110010010111",
452=>"0001010111000101",
453=>"1111000111111111",
454=>"1011010101011101",
455=>"1111101110100011",
456=>"0111100010001101",
457=>"0100101000100110",
458=>"1101001001010011",
459=>"1011101101001111",
460=>"1110111111101101",
461=>"0010001111001001",
462=>"0001001010100000",
463=>"1101110101000011",
464=>"1110010100100111",
465=>"0000011101100011",
466=>"0001010110100011",
467=>"0000000001011100",
468=>"1011110101001101",
469=>"1101110010001001",
470=>"0110010011101110",
471=>"0110010100110100",
472=>"1110100010000001",
473=>"1011011110111111",
474=>"1110000011010111",
475=>"0001101110111111",
476=>"0001110011110010",
477=>"1110011001010010",
478=>"1101110111111111",
479=>"0000000101010101",
480=>"0001001111111001",
481=>"0000101111000100",
482=>"1100101110011111",
483=>"1100011000010100",
484=>"0100100011100001",
485=>"0111100000111110",
486=>"0000010110000101",
487=>"1011011111010001",
488=>"1101001000111100",
489=>"0001000110000110",
490=>"0010010010010100",
491=>"1111001010001010",
492=>"1101100011101010",
493=>"1111100110011111",
494=>"0001000110001110",
495=>"0001001011010100",
496=>"1101110001010110",
497=>"1011011111100001",
498=>"0010011100101111",
499=>"0111111101010010",
500=>"0010010010000000",
501=>"1100000000100111",
502=>"1100011001000110",
503=>"0000001000111111",
504=>"0010100000010010",
505=>"0000000011110111",
506=>"1101011110110110",
507=>"1111000001000010",
508=>"0000111000010101",
509=>"0001010110010000",
510=>"1110111001000100",
511=>"1011010100011011",
512=>"0000001011110010",
513=>"0111101010110101",
514=>"0100001111100010",
515=>"1100111000110010",
516=>"1011110010101011",
517=>"1111001110110000",
518=>"0010010110100011",
519=>"0000111100010011",
520=>"1101101110001011",
521=>"1110011011111000",
522=>"0000100010000111",
523=>"0001011001011010",
524=>"1111111001001101",
525=>"1011101100000011",
526=>"1110001110101000",
527=>"0110101001100011",
528=>"0101111111001000",
529=>"1110001111110011",
530=>"1011011101001110",
531=>"1110010000111011",
532=>"0001110111100011",
533=>"0001110010111001",
534=>"1110010101000100",
535=>"1101111000000111",
536=>"0000000110001010",
537=>"0001001111000011",
538=>"0000101110011100",
539=>"1100100110100011",
540=>"1100011010011101",
541=>"0100101000100011",
542=>"0111011011011100",
543=>"0000010000010011",
544=>"1011100000011000",
545=>"1101001100111101",
546=>"0001000100011001",
547=>"0010010001111110",
548=>"1111001000111010",
549=>"1101100011010001",
550=>"1111101001001011",
551=>"0001000101011010",
552=>"0001001000001001",
553=>"1101101101011111",
554=>"1011100100000000",
555=>"0010100001101000",
556=>"0111111011101111",
557=>"0010001011010000",
558=>"1011111100111110",
559=>"1100011011011110",
560=>"0000001110101110",
561=>"0010011110111111",
562=>"0000000011110010",
563=>"1101011110101100",
564=>"1111000011101111",
565=>"0000111000111010",
566=>"0001010101010101",
567=>"1110110100011111",
568=>"1011010100100001",
569=>"0000010011001001",
570=>"0111101110001111",
571=>"0100001000110010",
572=>"1100110110010000",
573=>"1011110110010101",
574=>"1111010010100101",
575=>"0010010111100100",
576=>"0000111001101111",
577=>"1101101011010111",
578=>"1110011101101001",
579=>"0000100001011111",
580=>"0001011000010100",
581=>"1111110100001101",
582=>"1011101001010001",
583=>"1110010011111011",
584=>"0110101101111100",
585=>"0101111011100100",
586=>"1110001000110100",
587=>"1011011101101110",
588=>"1110010100101001",
589=>"0001111010111010",
590=>"0001101001001111",
591=>"1110001101011100",
592=>"1101111101000110",
593=>"0000001101100000",
594=>"0001001111000010",
595=>"0000100101011101",
596=>"1100011001110110",
597=>"1100101100111010",
598=>"0101000101111100",
599=>"0111001111100011",
600=>"1111110100110101",
601=>"1011011100110101",
602=>"1101011011011110",
603=>"0001001110010111",
604=>"0010001110011110",
605=>"1110111101110000",
606=>"1101101000101000",
607=>"1111101111010011",
608=>"0001000111100000",
609=>"0001000100110001",
610=>"1101011111001110",
611=>"1011101100100011",
612=>"0011000010001000",
613=>"0111111000100110",
614=>"0001110000001111",
615=>"1011110101010011",
616=>"1100100110001010",
617=>"0000011011010011",
618=>"0010011100110100",
619=>"1111110100011101",
620=>"1101011110110110",
621=>"1111001010110011",
622=>"0000111101000000",
623=>"0001010100000000",
624=>"1110100100100111",
625=>"1011010001001000",
626=>"0000110100010000",
627=>"0111110011010110",
628=>"0011110001101010",
629=>"1100100110110001",
630=>"1011111100011111",
631=>"1111100001001000",
632=>"0010010111000011",
633=>"0000101110001011",
634=>"1101100101100110",
635=>"1110101001001000",
636=>"0000100110010000",
637=>"0001011001101010",
638=>"1111100110001001",
639=>"1011011111010000",
640=>"1110011100111101",
641=>"0110110010101001",
642=>"0101110111001111",
643=>"1110000010111110",
644=>"1011011101111000",
645=>"1110010111110000",
646=>"0001111111110101",
647=>"0001100101101101",
648=>"1110001011001000",
649=>"1110000000010010",
650=>"0000001111011110",
651=>"0001010100001111",
652=>"0000100011000010",
653=>"1100010110001111",
654=>"1100110010000011",
655=>"0101001101110000",
656=>"0111001001110110",
657=>"1111101101010000",
658=>"1011011110110111",
659=>"1101011011000101",
660=>"0001010010101100",
661=>"0010001101011111",
662=>"1110111000010010",
663=>"1101100111011010",
664=>"1111110000100000",
665=>"0001001011010001",
666=>"0001000001011101",
667=>"1101011011111000",
668=>"1011101101100110",
669=>"0011001000100000",
670=>"0111110111111101",
671=>"0001100111011001",
672=>"1011110001110011",
673=>"1100100111010100",
674=>"0000011111110011",
675=>"0010011110000010",
676=>"1111110000001100",
677=>"1101011110100010",
678=>"1111001100010000",
679=>"0000111011001110",
680=>"0001010101101000",
681=>"1110100011111101",
682=>"1011010011110100",
683=>"0000111110010110",
684=>"0111110110000000",
685=>"0011101000001100",
686=>"1100100010111111",
687=>"1011111101110100",
688=>"1111100010011001",
689=>"0010011010001011",
690=>"0000100111101111",
691=>"1101101000000001",
692=>"1110101010111010",
693=>"0000101001101010",
694=>"0001011000101111",
695=>"1111100011001111",
696=>"1011011100111101",
697=>"1110110101001001",
698=>"0111000100001101",
699=>"0101011111011111",
700=>"1101101101101110",
701=>"1011100100000000",
702=>"1110100100110110",
703=>"0010000101101011",
704=>"0001100001011011",
705=>"1110000010011100",
706=>"1110000111100001",
707=>"0000010011110010",
708=>"0001010100100000",
709=>"0000010111111010",
710=>"1100001011110111",
711=>"1101000100011011",
712=>"0101100111111011",
713=>"0110111001001000",
714=>"1111010010101111",
715=>"1011011011110110",
716=>"1101101000100011",
717=>"0001011100101000",
718=>"0010000110001010",
719=>"1110101111110001",
720=>"1101101011100011",
721=>"1111110110111101",
722=>"0001001010110100",
723=>"0000111011100111",
724=>"1101001010011110",
725=>"1011111001010010",
726=>"0011100110011001",
727=>"0111110011000101",
728=>"0001001001000111",
729=>"1011101100010101",
730=>"1100110100100011",
731=>"0000101001110000",
732=>"0010011000100110",
733=>"1111100011011110",
734=>"1101100000100011",
735=>"1111010111000010",
736=>"0000111110100000",
737=>"0001010001011010",
738=>"1110010010111100",
739=>"1011010111111110",
740=>"0001011100001000",
741=>"0111111101011000",
742=>"0011001100101111",
743=>"1100010100101010",
744=>"1100000100000001",
745=>"1111110011100001",
746=>"0010011100100100",
747=>"0000100110101101",
748=>"1101100101110010",
749=>"1110101011001001",
750=>"0000101010101001",
751=>"0001010101110011",
752=>"1111100001101100",
753=>"1011011011110000",
754=>"1110111101101101",
755=>"0111000111111011",
756=>"0101011001010110",
757=>"1101101001000010",
758=>"1011100101100111",
759=>"1110101001000111",
760=>"0010000011111101",
761=>"0001011101110010",
762=>"1110000001101110",
763=>"1110001010001101",
764=>"0000010100110110",
765=>"0001010100101101",
766=>"0000010110110000",
767=>"1100001001000001",
768=>"1101001100100001",
769=>"0101101011100111",
770=>"0110110101100000",
771=>"1111001111011010",
772=>"1011011100011111",
773=>"1101101100101111",
774=>"0001100000001001",
775=>"0010000011000001",
776=>"1110101011111000",
777=>"1101101100101100",
778=>"1111111001010000",
779=>"0001001110011010",
780=>"0000111010000101",
781=>"1101000101110001",
782=>"1011111011000101",
783=>"0011101111110010",
784=>"0111101110111000",
785=>"0001001001100000",
786=>"1011101000000011",
787=>"1100110111111110",
788=>"0000101101011010",
789=>"0010011001010001",
790=>"1111011111111101",
791=>"1101011110011011",
792=>"1111011000111111",
793=>"0000111101001010",
794=>"0001010010000100",
795=>"1110001100100010",
796=>"1011010101000111",
797=>"0001100011000100",
798=>"0111111010110010",
799=>"0011000101111101",
800=>"1100010010111010",
801=>"1100001000101100",
802=>"1111110011001101",
803=>"0010011011101000",
804=>"0000011011110000",
805=>"1101100010011011",
806=>"1110110100101111",
807=>"0000101111111111",
808=>"0001010111100110",
809=>"1111010001001000",
810=>"1011011001110001",
811=>"1111011001011101",
812=>"0111010101001101",
813=>"0100111101101000",
814=>"1101010110110101",
815=>"1011101001011111",
816=>"1110110110011111",
817=>"0010001100100010",
818=>"0001010011001011",
819=>"1101111010000100",
820=>"1110001110101101",
821=>"0000011100010011",
822=>"0001010110101101",
823=>"0000001001101100",
824=>"1011111110001100",
825=>"1101100000100111",
826=>"0110000011101001",
827=>"0110100011101100",
828=>"1110110101101001",
829=>"1011011101100001",
830=>"1101111001101000",
831=>"0001101011111000",
832=>"0001111100011101",
833=>"1110011111010000",
834=>"1101110000110110",
835=>"1111111101101010",
836=>"0001001101000100",
837=>"0000110101100100",
838=>"1100110111011010",
839=>"1100001011110001",
840=>"0100001101010000",
841=>"0111101000011100",
842=>"0000101001111100",
843=>"1011100011001101",
844=>"1101000000110000",
845=>"0000111011010011",
846=>"0010010100101111",
847=>"1111010100111000",
848=>"1101011111110100",
849=>"1111100000110101",
850=>"0001000000010111",
851=>"0001001011110001",
852=>"1110000000011001",
853=>"1011010101110010",
854=>"0001101011001011",
855=>"0111111110000000",
856=>"0010111110110001",
857=>"1100001101111011",
858=>"1100001011111111",
859=>"1111110110101011",
860=>"0010100000001101",
861=>"0000011001100011",
862=>"1101100010010001",
863=>"1110110110010000",
864=>"0000110000010000",
865=>"0001010111101001",
866=>"1111001110110111",
867=>"1011010111011111",
868=>"1111011111101110",
869=>"0111011100010010",
870=>"0100110101001101",
871=>"1101010010000010",
872=>"1011101010010111",
873=>"1110111001000111",
874=>"0010001100010101",
875=>"0001010000001001",
876=>"1101111000001100",
877=>"1110010001000001",
878=>"0000011010111011",
879=>"0001010110001100",
880=>"0000000110110111",
881=>"1011111010011011",
882=>"1101100110001111",
883=>"0110001000111111",
884=>"0110011110101000",
885=>"1110101101011110",
886=>"1011011110001010",
887=>"1101111101000111",
888=>"0001101010011110",
889=>"0001111000000001",
890=>"1110011101111110",
891=>"1101110101011000",
892=>"0000000010000011",
893=>"0001001111000000",
894=>"0000110010101001",
895=>"1100110101110001",
896=>"1100010000010011",
897=>"0100010101100110",
898=>"0111100110011001",
899=>"0000100011100101",
900=>"1011100001001010",
901=>"1101000011001010",
902=>"0001000000001111",
903=>"0010010100110001",
904=>"1111001111111010",
905=>"1101100010101000",
906=>"1111100010100010",
907=>"0001000100111111",
908=>"0001001101001011",
909=>"1101111001011101",
910=>"1011011011110101",
911=>"0010001101011100",
912=>"0111111101100100",
913=>"0010100000001001",
914=>"1100000101010010",
915=>"1100010100101101",
916=>"0000000010010000",
917=>"0010100000011001",
918=>"0000001010000100",
919=>"1101011111110000",
920=>"1110111100110000",
921=>"0000110110101010",
922=>"0001010110110001",
923=>"1111000000100001",
924=>"1011010101001101",
925=>"1111111101000101",
926=>"0111100101100111",
927=>"0100011100111001",
928=>"1101000000100010",
929=>"1011101111110010",
930=>"1111000111101000",
931=>"0010010100101100",
932=>"0001000001110101",
933=>"1101110001010000",
934=>"1110010111101111",
935=>"0000100000000011",
936=>"0001011000101000",
937=>"1111111111100101",
938=>"1011110000001001",
939=>"1110000010011101",
940=>"0110011111010010",
941=>"0110001010010001",
942=>"1110011001111101",
943=>"1011011100111101",
944=>"1110001001001011",
945=>"0001110101010111",
946=>"0001101111010000",
947=>"1110010011000101",
948=>"1101111011110011",
949=>"0000001000001001",
950=>"0001010000111001",
951=>"0000101011000011",
952=>"1100100011001110",
953=>"1100011110001001",
954=>"0100110001001101",
955=>"0111011010010011",
956=>"0000000111111111",
957=>"1011011110100010",
958=>"1101010001000111",
959=>"0001000000001110",
960=>"0010010011111110",
961=>"1111001110111100",
962=>"1101100001111100",
963=>"1111100101011010",
964=>"0001000100000101",
965=>"0001001010001110",
966=>"1101110101010100",
967=>"1011100000010100",
968=>"0010010010010001",
969=>"0111111100011010",
970=>"0010011001001110",
971=>"1100000001101110",
972=>"1100010110101100",
973=>"0000001000010001",
974=>"0010011111000001",
975=>"0000001010000111",
976=>"1101011111011000",
977=>"1110111111101000",
978=>"0000110111000110",
979=>"0001010110001000",
980=>"1110111011101111",
981=>"1011010101010101",
982=>"0000000100000101",
983=>"0111101001100010",
984=>"0100010110000000",
985=>"1100111110000001",
986=>"1011110011000110",
987=>"1111001011110011",
988=>"0010010101011111",
989=>"0000111111101011",
990=>"1101101101111111",
991=>"1110011001110100",
992=>"0000011111001001",
993=>"0001010111111100",
994=>"1111111010010010",
995=>"1011101101100100",
996=>"1110000111001100",
997=>"0110100100010101",
998=>"0110000110010101",
999=>"1110010011100110",
1000=>"1011011100011011",
1001=>"1110001110000000",
1002=>"0001110111000010",
1003=>"0001101101110001",
1004=>"1110010001111100",
1005=>"1101111001111110",
1006=>"0000001010100011",
1007=>"0001001110001011",
1008=>"0000101001100110",
1009=>"1100100000110000",
1010=>"1100100011101001",
1011=>"0100111000110000",
1012=>"0111010110010001",
1013=>"0000000001111001",
1014=>"1011011101110111",
1015=>"1101010101100100",
1016=>"0001001000111101",
1017=>"0010010001001010",
1018=>"1111000011100000",
1019=>"1101100110111111",
1020=>"1111101011101101",
1021=>"0001000110001110",
1022=>"0001000111001001",
1023=>"1101100111000110");
  
  rom1 <= (
0=>"1011100111110001",
1=>"0010110011000000",
2=>"0111111010011000",
3=>"0001111110001101",
4=>"1011111001010100",
5=>"1100100001001110",
6=>"0000010100111001",
7=>"0010011101100000",
8=>"1111111010100111",
9=>"1101011111001100",
10=>"1111000110100111",
11=>"0000111011011001",
12=>"0001010100111100",
13=>"1110101100010100",
14=>"1011010000110000",
15=>"0000100101000110",
16=>"0111101111101100",
17=>"0011111111001101",
18=>"1100101101111100",
19=>"1011111000111000",
20=>"1111011010010101",
21=>"0010010101100111",
22=>"0000110011111110",
23=>"1101101000000101",
24=>"1110100100110010",
25=>"0000100100100100",
26=>"0001011000111010",
27=>"1111101101010100",
28=>"1011100010101000",
29=>"1110100000110100",
30=>"0110110101101101",
31=>"0101101111001010",
32=>"1101111111100001",
33=>"1011100000011101",
34=>"1110011010110111",
35=>"0001111101001100",
36=>"0001100110010011",
37=>"1110001000100111",
38=>"1110000010000001",
39=>"0000010000111111",
40=>"0001010010111000",
41=>"0000011111010000",
42=>"1100011011110100",
43=>"1100101001000000",
44=>"0101000000011101",
45=>"0111010001001001",
46=>"1111111001111000",
47=>"1011011111111111",
48=>"1101010101000011",
49=>"0001001101010011",
50=>"0010010000010101",
51=>"1110111110000101",
52=>"1101100101100101",
53=>"1111101100111001",
54=>"0001001001111111",
55=>"0001000100000101",
56=>"1101100011100010",
57=>"1011101000110100",
58=>"0010111001001100",
59=>"0111111010001101",
60=>"0001110101010000",
61=>"1011110101101111",
62=>"1100100010001001",
63=>"0000011001100000",
64=>"0010011110101111",
65=>"1111110110100011",
66=>"1101011110100011",
67=>"1111001000010101",
68=>"0000111001011100",
69=>"0001010110101001",
70=>"1110101011100110",
71=>"1011010011011000",
72=>"0000101110111101",
73=>"0111110010111011",
74=>"0011110101101010",
75=>"1100101010000011",
76=>"1011111010000011",
77=>"1111011011101100",
78=>"0010011000101011",
79=>"0000101101111000",
80=>"1101101001111011",
81=>"1110100111000011",
82=>"0000100111011101",
83=>"0001011000101100",
84=>"1111101001110000",
85=>"1011100000011010",
86=>"1110100111011111",
87=>"0110111011111001",
88=>"0101101011000011",
89=>"1101110111110011",
90=>"1011100001111111",
91=>"1110011110010010",
92=>"0010000010000000",
93=>"0001100110100100",
94=>"1110000110011010",
95=>"1110000100001101",
96=>"0000010000111011",
97=>"0001010011110101",
98=>"0000011100100101",
99=>"1100010010001011",
100=>"1100111010000111",
101=>"0101011011100010",
102=>"0111000001010010",
103=>"1111011111000100",
104=>"1011011100010000",
105=>"1101100010011001",
106=>"0001010111100001",
107=>"0010001001011011",
108=>"1110110101001111",
109=>"1101101001100001",
110=>"1111110011011101",
111=>"0001001001101011",
112=>"0000111110100000",
113=>"1101010010001001",
114=>"1011110011010101",
115=>"0011010111100001",
116=>"0111110110010111",
117=>"0001010111000011",
118=>"1011101111010100",
119=>"1100101111011001",
120=>"0000100011100011",
121=>"0010011001111010",
122=>"1111101001100000",
123=>"1101100000010100",
124=>"1111010010111101",
125=>"0000111101000111",
126=>"0001010010100001",
127=>"1110011010111001",
128=>"1011010110010100",
129=>"0001001100111011",
130=>"0111111011000010",
131=>"0011011010111100",
132=>"1100011010100111",
133=>"1100000000011010",
134=>"1111101100000100",
135=>"0010011100100011",
136=>"0000100001110010",
137=>"1101100110000111",
138=>"1110101101110000",
139=>"0000101101111100",
140=>"0001011001100101",
141=>"1111011101000111",
142=>"1011011010011010",
143=>"1111000101100111",
144=>"0111001100101101",
145=>"0101010000001000",
146=>"1101100100110000",
147=>"1011101000001011",
148=>"1110100100100101",
149=>"0001111111110111",
150=>"0001100011001111",
151=>"1110000101010110",
152=>"1110000111000010",
153=>"0000010001111010",
154=>"0001010100001000",
155=>"0000011011011100",
156=>"1100001111010000",
157=>"1101000001111101",
158=>"0101011111100100",
159=>"0110111101101010",
160=>"1111011011101111",
161=>"1011011100101101",
162=>"1101100110100101",
163=>"0001011011000111",
164=>"0010000110011111",
165=>"1110110001001100",
166=>"1101101010100111",
167=>"1111110101101001",
168=>"0001001101010110",
169=>"0000111101000111",
170=>"1101001101011100",
171=>"1011110100110001",
172=>"0011100001000100",
173=>"0111110010010111",
174=>"0001010111010010",
175=>"1011101011001100",
176=>"1100110010011101",
177=>"0000100111011111",
178=>"0010011010011111",
179=>"1111100110010010",
180=>"1101011101110011",
181=>"1111010101001010",
182=>"0000111011100100",
183=>"0001010011011011",
184=>"1110010100011100",
185=>"1011010011010110",
186=>"0001010011100111",
187=>"0111111001000011",
188=>"0011010011110000",
189=>"1100011001000101",
190=>"1100000100100001",
191=>"1111101100100110",
192=>"0010011010101100",
193=>"0000100001111101",
194=>"1101100011111111",
195=>"1110110000101000",
196=>"0000101110000011",
197=>"0001010111110001",
198=>"1111011000000010",
199=>"1011011100000110",
200=>"1111001011010110",
201=>"0111001110001101",
202=>"0101001001111110",
203=>"1101011111111100",
204=>"1011100111000101",
205=>"1110101111101100",
206=>"0010001001100111",
207=>"0001011000011101",
208=>"1101111101101101",
209=>"1110001011000010",
210=>"0000011001101011",
211=>"0001010110001011",
212=>"0000001110111101",
213=>"1100000011101011",
214=>"1101010101011111",
215=>"0101111000000100",
216=>"0110101101000010",
217=>"1111000001010001",
218=>"1011011101010111",
219=>"1101110011001011",
220=>"0001100111010001",
221=>"0010000000010001",
222=>"1110100100011111",
223=>"1101101110001110",
224=>"1111111010100000",
225=>"0001001011110001",
226=>"0000111001000111",
227=>"1100111110101100",
228=>"1100000100101010",
229=>"0011111110110001",
230=>"0111101101010000",
231=>"0000110111011001",
232=>"1011100101110001",
233=>"1100111010111010",
234=>"0000110101101001",
235=>"0010010110010111",
236=>"1111011011001010",
237=>"1101011110101100",
238=>"1111011101010010",
239=>"0000111110100010",
240=>"0001001110001100",
241=>"1110000110001000",
242=>"1011010111010111",
243=>"0001110100111101",
244=>"0111111101100101",
245=>"0010110111111001",
246=>"1100001010110100",
247=>"1100001111100100",
248=>"1111111001101000",
249=>"0010011101000101",
250=>"0000010110011010",
251=>"1101100010111000",
252=>"1110111000111110",
253=>"0000110000110010",
254=>"0001010111100011",
255=>"1111010101111010",
256=>"1011011001101110",
257=>"1111010001010110",
258=>"0111010101100110",
259=>"0101000001110001",
260=>"1101011010111010",
261=>"1011100111111000",
262=>"1110110010010101",
263=>"0010001001011111",
264=>"0001010101011110",
265=>"1101111011101101",
266=>"1110001101010110",
267=>"0000011000011000",
268=>"0001010101100110",
269=>"0000001100010010",
270=>"1011111111110001",
271=>"1101011010111001",
272=>"0101111101101000",
273=>"0110101000001100",
274=>"1110111001000000",
275=>"1011011101110000",
276=>"1101110110101111",
277=>"0001100101111110",
278=>"0001111011110111",
279=>"1110100011000000",
280=>"1101110010101111",
281=>"1111111110111001",
282=>"0001001101111000",
283=>"0000110110001110",
284=>"1100111101000000",
285=>"1100001000111100",
286=>"0100000111010000",
287=>"0111101011011101",
288=>"0000110001000100",
289=>"1011100011100010",
290=>"1100111101010100",
291=>"0000111010011100",
292=>"0010010110110010",
293=>"1111010101111011",
294=>"1101100001100101",
295=>"1111011110110000",
296=>"0001000011100000",
297=>"0001001111000011",
298=>"1110000001010111",
299=>"1011011000110110",
300=>"0001111101111001",
301=>"0111111101011110",
302=>"0010101110000100",
303=>"1100001010100000",
304=>"1100010000010000",
305=>"1111111011101010",
306=>"0010100000000011",
307=>"0000010000011110",
308=>"1101100000101010",
309=>"1110111000101101",
310=>"0000110100101101",
311=>"0001010111011000",
312=>"1111000111100111",
313=>"1011010110101011",
314=>"1111101110010010",
315=>"0111100000000011",
316=>"0100101001110100",
317=>"1101001000110111",
318=>"1011101100110100",
319=>"1111000000110011",
320=>"0010010010010100",
321=>"0001000111100010",
322=>"1101110100001101",
323=>"1110010100000000",
324=>"0000011101100011",
325=>"0001011000001010",
326=>"0000000101010111",
327=>"1011110100111111",
328=>"1101110110001011",
329=>"0110010101000100",
330=>"0110010100011101",
331=>"1110100101000110",
332=>"1011011100000110",
333=>"1110000010100111",
334=>"0001110001001010",
335=>"0001110011100111",
336=>"1110010111101110",
337=>"1101111000111000",
338=>"0000000101001010",
339=>"0001001111110101",
340=>"0000101111000101",
341=>"1100101010010000",
342=>"1100010101101101",
343=>"0100100011011001",
344=>"0111100000011010",
345=>"0000010101001010",
346=>"1011100000001101",
347=>"1101001011001001",
348=>"0001000010110001",
349=>"0010010111010011",
350=>"1111001011100001",
351=>"1101100011101000",
352=>"1111100101111110",
353=>"0001000100111000",
354=>"0001001001010000",
355=>"1101110010101001",
356=>"1011011111100011",
357=>"0010011011110111",
358=>"0111111110010111",
359=>"0010001111010010",
360=>"1011111111111111",
361=>"1100010101000110",
362=>"0000000000111110",
363=>"0010011111001111",
364=>"0000010000001010",
365=>"1101100000100000",
366=>"1110111011010100",
367=>"0000110101011001",
368=>"0001010110101001",
369=>"1111000011000010",
370=>"1011010110011011",
371=>"1111110101010110",
372=>"0111100100001001",
373=>"0100100011001010",
374=>"1101000110000001",
375=>"1011110000001100",
376=>"1111000100111001",
377=>"0010010011010011",
378=>"0001000101011000",
379=>"1101110000111100",
380=>"1110010101111100",
381=>"0000011100110100",
382=>"0001010111011001",
383=>"0000000000010010",
384=>"1011110010000110",
385=>"1101111010111000",
386=>"0110011010001001",
387=>"0110010000110101",
388=>"1110011110100010",
389=>"1011011011011110",
390=>"1110000111010001",
391=>"0001110011000101",
392=>"0001110010000000",
393=>"1110010110101110",
394=>"1101110110111000",
395=>"0000000111101000",
396=>"0001001101001011",
397=>"0000101101101000",
398=>"1100100111101101",
399=>"1100011010111100",
400=>"0100101011001010",
401=>"0111011100101000",
402=>"0000001111000000",
403=>"1011011111010100",
404=>"1101001111101000",
405=>"0001000011100010",
406=>"0010010011011111",
407=>"1111001001011111",
408=>"1101100101011000",
409=>"1111101000001011",
410=>"0001000100110010",
411=>"0001001001011110",
412=>"1101101110111000",
413=>"1011100011101001",
414=>"0010100011100111",
415=>"0111111011101111",
416=>"0010001100000100",
417=>"1011111101110010",
418=>"1100011100010000",
419=>"0000001110100100",
420=>"0010011101110010",
421=>"0000000000111110",
422=>"1101011111100100",
423=>"1111000010100110",
424=>"0000111001100011",
425=>"0001010101111010",
426=>"1110110011110000",
427=>"1011010001000011",
428=>"0000010101110101",
429=>"0111101011101100",
430=>"0100001100010111",
431=>"1100110101101100",
432=>"1011110101001101",
433=>"1111010011110010",
434=>"0010010011101010",
435=>"0000111010000001",
436=>"1101101010011010",
437=>"1110100000111001",
438=>"0000100010010100",
439=>"0001011000101000",
440=>"1111110011101000",
441=>"1011100110100110",
442=>"1110010011101010",
443=>"0110101100101100",
444=>"0101111010001001",
445=>"1110001010000010",
446=>"1011011110110111",
447=>"1110010100010011",
448=>"0001111001010111",
449=>"0001101011000100",
450=>"1110001100111000",
451=>"1101111110110110",
452=>"0000001101111110",
453=>"0001010010010100",
454=>"0000100010110100",
455=>"1100011011010011",
456=>"1100101110010110",
457=>"0101000100100110",
458=>"0111001100111001",
459=>"1111110011011111",
460=>"1011011101011111",
461=>"1101011001110110",
462=>"0001010001001011",
463=>"0010001110100111",
464=>"1110111110000110",
465=>"1101100110000000",
466=>"1111101111110100",
467=>"0001001001100001",
468=>"0001000110011011",
469=>"1101101011010001",
470=>"1011100100100001",
471=>"0010101001110010",
472=>"0111111011111000",
473=>"0010000011001010",
474=>"1011111010000001",
475=>"1100011101001000",
476=>"0000010011000101",
477=>"0010011111001111",
478=>"1111111100111000",
479=>"1101011110110100",
480=>"1111000100010101",
481=>"0000110111101010",
482=>"0001010111011111",
483=>"1110110011001011",
484=>"1011010011010111",
485=>"0000011111101111",
486=>"0111101111001011",
487=>"0100000011000011",
488=>"1100110001011011",
489=>"1011110110100000",
490=>"1111010100111100",
491=>"0010010110111111",
492=>"0000110011111000",
493=>"1101101100000111",
494=>"1110100011001010",
495=>"0000100101010000",
496=>"0001011000011111",
497=>"1111110000001001",
498=>"1011100100001011",
499=>"1110011010001100",
500=>"0110110011000010",
501=>"0101110110010111",
502=>"1110000010000111",
503=>"1011100000010000",
504=>"1110010111101011",
505=>"0001111110001101",
506=>"0001101011011110",
507=>"1110001010101000",
508=>"1110000000111011",
509=>"0000001110000110",
510=>"0001010011000000",
511=>"0000100001001001",
512=>"1100011000101000",
513=>"1100110000010101",
514=>"0101001110101010",
515=>"0111001001000101",
516=>"1111101011100010",
517=>"1011011101000011",
518=>"1101011100001101",
519=>"0001010010011000",
520=>"0010001100010111",
521=>"1110111010111100",
522=>"1101100111100011",
523=>"1111101111111110",
524=>"0001001000011001",
525=>"0001000001010100",
526=>"1101011001110000",
527=>"1011101101111111",
528=>"0011001000010110",
529=>"0111111001001101",
530=>"0001100100111001",
531=>"1011110010110001",
532=>"1100101010001101",
533=>"0000011101011010",
534=>"0010011010110110",
535=>"1111101111110000",
536=>"1101100000000101",
537=>"1111001111000011",
538=>"0000111011011101",
539=>"0001010011101111",
540=>"1110100010100001",
541=>"1011010101011010",
542=>"0000111101100000",
543=>"0111111000011010",
544=>"0011101000101010",
545=>"1100100001010110",
546=>"1011111100011010",
547=>"1111100101010011",
548=>"0010011011011100",
549=>"0000100111111001",
550=>"1101100111111011",
551=>"1110101001110010",
552=>"0000101011110010",
553=>"0001011001101010",
554=>"1111100011110010",
555=>"1011011101011111",
556=>"1110110111100110",
557=>"0111000101001000",
558=>"0101011011110111",
559=>"1101101110101000",
560=>"1011100101011011",
561=>"1110100010110011",
562=>"0010000101010100",
563=>"0001011110101111",
564=>"1110000001100110",
565=>"1110000101111010",
566=>"0000010101000001",
567=>"0001010110000001",
568=>"0000010111001100",
569=>"1100001100101010",
570=>"1101000101001111",
571=>"0101100101101001",
572=>"0110111001011000",
573=>"1111010011010100",
574=>"1011011001100111",
575=>"1101100000110010",
576=>"0001010101110111",
577=>"0010001001101111",
578=>"1110110110101010",
579=>"1101101000101011",
580=>"1111110010000010",
581=>"0001001100001011",
582=>"0000111111111111",
583=>"1101010101001010",
584=>"1011101111000000",
585=>"0011010010000111",
586=>"0111110101010110",
587=>"0001100101000100",
588=>"1011101110101110",
589=>"1100101100111111",
590=>"0000100001100001",
591=>"0010011011011011",
592=>"1111101100101011",
593=>"1101011101011001",
594=>"1111010001010011",
595=>"0000111001111011",
596=>"0001010100101010",
597=>"1110011100010010",
598=>"1011010010000110",
599=>"0001000100001011",
600=>"0111110110101110",
601=>"0011100001011011",
602=>"1100011111101000",
603=>"1100000000011111",
604=>"1111100101111101",
605=>"0010011001100001",
606=>"0000101000000111",
607=>"1101100101101110",
608=>"1110101100100100",
609=>"0000101100000010",
610=>"0001010111110111",
611=>"1111011110110001",
612=>"1011011110110111",
613=>"1110111101011101",
614=>"0111000110101101",
615=>"0101010110000001",
616=>"1101101001011001",
617=>"1011100100110110",
618=>"1110101000111101",
619=>"0010000110011100",
620=>"0001011101101001",
621=>"1110000001100000",
622=>"1110000111011111",
623=>"0000010110111100",
624=>"0001010101100101",
625=>"0000010100000001",
626=>"1100001001011101",
627=>"1101001010101101",
628=>"0101101100001001",
629=>"0110110101111001",
630=>"1111001101001100",
631=>"1011011101011100",
632=>"1101101100110011",
633=>"0001100010011101",
634=>"0010000011111011",
635=>"1110101001110100",
636=>"1101101011110011",
637=>"1111110111001110",
638=>"0001001010100001",
639=>"0000111100011001",
640=>"1101000110001011",
641=>"1011111101111110",
642=>"0011110000001000",
643=>"0111110001011101",
644=>"0001000101000011",
645=>"1011101000100100",
646=>"1100110101010010",
647=>"0000101111101110",
648=>"0010010111111100",
649=>"1111100001010100",
650=>"1101011110000000",
651=>"1111011001010111",
652=>"0000111101001001",
653=>"0001001111100111",
654=>"1110001110000110",
655=>"1011010101000101",
656=>"0001100101011101",
657=>"0111111100011100",
658=>"0011000101110111",
659=>"1100010000100110",
660=>"1100001011001001",
661=>"1111110011001100",
662=>"0010011100010000",
663=>"0000011100110000",
664=>"1101100100000010",
665=>"1110110101001010",
666=>"0000101110100001",
667=>"0001011000011111",
668=>"1111010010110110",
669=>"1011011001101011",
670=>"1111011010101010",
671=>"0111010110001111",
672=>"0100111101101010",
673=>"1101011000000010",
674=>"1011101010000111",
675=>"1110110110110100",
676=>"0010001011110100",
677=>"0001010000011101",
678=>"1101111001101110",
679=>"1110001110101100",
680=>"0000011011101110",
681=>"0001010111110101",
682=>"0000010000101111",
683=>"1100000101110111",
684=>"1101001111100100",
685=>"0101110010001100",
686=>"0110110001000101",
687=>"1111000101000001",
688=>"1011011101011010",
689=>"1101110000100111",
690=>"0001100001001000",
691=>"0001111111101100",
692=>"1110101000000001",
693=>"1101110000011000",
694=>"1111111011100001",
695=>"0001001100110101",
696=>"0000111001011110",
697=>"1101000100011110",
698=>"1100000001111101",
699=>"0011111000110011",
700=>"0111101111110111",
701=>"0000111110110000",
702=>"1011100110000111",
703=>"1100110111101010",
704=>"0000110100011100",
705=>"0010011000101001",
706=>"1111011011111100",
707=>"1101100000110100",
708=>"1111011010110100",
709=>"0001000010000100",
710=>"0001010000101011",
711=>"1110001001010101",
712=>"1011010110010011",
713=>"0001101110011000",
714=>"0111111100101110",
715=>"0010111100000000",
716=>"1100010000000000",
717=>"1100001100000000",
718=>"1111110100111110",
719=>"0010011111100000",
720=>"0000010110110011",
721=>"1101100001110101",
722=>"1110110100100110",
723=>"0000110010110000",
724=>"0001010111110100",
725=>"1111001110101001",
726=>"1011011000100001",
727=>"1111011111101111",
728=>"0111011001111010",
729=>"0100110110100011",
730=>"1101010001011101",
731=>"1011101010000110",
732=>"1110111001111100",
733=>"0010001111110000",
734=>"0001001101000110",
735=>"1101110111011010",
736=>"1110010000010011",
737=>"0000011011000010",
738=>"0001010111100100",
739=>"0000001010111111",
740=>"1011111010000110",
741=>"1101101010010010",
742=>"0110001010011001",
743=>"0110011110010000",
744=>"1110110000011110",
745=>"1011011011100001",
746=>"1101111100000101",
747=>"0001101100110011",
748=>"0001110111110010",
749=>"1110011100100001",
750=>"1101110110000110",
751=>"0000000010000100",
752=>"0001001110110000",
753=>"0000110010111001",
754=>"1100110001011101",
755=>"1100001101101101",
756=>"0100010101010110",
757=>"0111100101111101",
758=>"0000100010100100",
759=>"1011100010000110",
760=>"1101000101011001",
761=>"0000111101000000",
762=>"0010011001011100",
763=>"1111010001100111",
764=>"1101100010011001",
765=>"1111100010001101",
766=>"0001000011100000",
767=>"0001001011001110",
768=>"1101111010100011",
769=>"1011011100000100",
770=>"0010001100011010",
771=>"0111111110101101",
772=>"0010011101100110",
773=>"1100000100001011",
774=>"1100010011111000",
775=>"0000000100000101",
776=>"0010011101100110",
777=>"0000001100111010",
778=>"1101011111111111",
779=>"1110111101011001",
780=>"0000110011010111",
781=>"0001010110100011",
782=>"1110111110011100",
783=>"1011010101001010",
784=>"1111111100101010",
785=>"0111100111001000",
786=>"0100011011001001",
787=>"1101000000001111",
788=>"1011101110100000",
789=>"1110111101100100",
790=>"0010010001000111",
791=>"0001001010110110",
792=>"1101110100001101",
793=>"1110010010000011",
794=>"0000011010011110",
795=>"0001010110101111",
796=>"0000000110000101",
797=>"1011110110111101",
798=>"1101101110111010",
799=>"0110001111100010",
800=>"0110011010111100",
801=>"1110101001110000",
802=>"1011011010110001",
803=>"1110000000101000",
804=>"0001101110111011",
805=>"0001110110000111",
806=>"1110011011100111",
807=>"1101110011111110",
808=>"0000000100100101",
809=>"0001001100001010",
810=>"0000110001011010",
811=>"1100101110111010",
812=>"1100010010101010",
813=>"0100011101010100",
814=>"0111100010011011",
815=>"0000011100010100",
816=>"1011100001000010",
817=>"1101001001110100",
818=>"0000111101111101",
819=>"0010010101100111",
820=>"1111001111100010",
821=>"1101100100000000",
822=>"1111100100100010",
823=>"0001000011010111",
824=>"0001001011100011",
825=>"1101110110101101",
826=>"1011011111111110",
827=>"0010010100001101",
828=>"0111111100011110",
829=>"0010011001111110",
830=>"1100000010100100",
831=>"1100010111011101",
832=>"0000001000001010",
833=>"0010011101110111",
834=>"0000000111010001",
835=>"1101100000001110",
836=>"1110111110100001",
837=>"0000110111101100",
838=>"0001010110101101",
839=>"1110111011000111",
840=>"1011010001110001",
841=>"0000000110110000",
842=>"0111100111000100",
843=>"0100011001011001",
844=>"1100111101101111",
845=>"1011110001101111",
846=>"1111001101001100",
847=>"0010010001100001",
848=>"0000111111111011",
849=>"1101101101000000",
850=>"1110011101000000",
851=>"0000100000000100",
852=>"0001011000001101",
853=>"1111111001110001",
854=>"1011101010111001",
855=>"1110000110110111",
856=>"0110100011001001",
857=>"0110000100110110",
858=>"1110010100110001",
859=>"1011011101100100",
860=>"1110001101101111",
861=>"0001110101011010",
862=>"0001101111100110",
863=>"1110010001011001",
864=>"1101111011101101",
865=>"0000001011000000",
866=>"0001010001011101",
867=>"0000100111000110",
868=>"1100100001111111",
869=>"1100100101010001",
870=>"0100110111010111",
871=>"0111010011101111",
872=>"0000000000011000",
873=>"1011011110101000",
874=>"1101010011110111",
875=>"0001001011101110",
876=>"0010010001010111",
877=>"1111000011110101",
878=>"1101100100011111",
879=>"1111101011111010",
880=>"0001001000110000",
881=>"0001000100101100",
882=>"1101100110100100",
883=>"1011100111001001",
884=>"0010110001110010",
885=>"0111111100001101",
886=>"0001111011101011",
887=>"1011111001101111",
888=>"1100100001010011",
889=>"0000010110100101",
890=>"0010011111001111",
891=>"1111111001100010",
892=>"1101011101001010",
893=>"1111000110011001",
894=>"0000110110000100",
895=>"0001011000010010",
896=>"1110111010100100",
897=>"1011010011111010",
898=>"0000010000100011",
899=>"0111101010111101",
900=>"0100010000001100",
901=>"1100111001001101",
902=>"1011110011000101",
903=>"1111001110001100",
904=>"0010010101000011",
905=>"0000111001110110",
906=>"1101101110011101",
907=>"1110011111010111",
908=>"0000100010111100",
909=>"0001011000001110",
910=>"1111110110010101",
911=>"1011101000010110",
912=>"1110001101001011",
913=>"0110101001101101",
914=>"0110000001010011",
915=>"1110001100110001",
916=>"1011011110101111",
917=>"1110010001001001",
918=>"0001111010001101",
919=>"0001110000001111",
920=>"1110001111000000",
921=>"1101111101110010",
922=>"0000001011001001",
923=>"0001010010001010",
924=>"0000100101011110",
925=>"1100011111010011",
926=>"1100100110111110",
927=>"0101000001011111",
928=>"0111010000010111",
929=>"1111111000001101",
930=>"1011011110000110",
931=>"1101010110001001",
932=>"0001001101000101",
933=>"0010001111000111",
934=>"1111000000101110",
935=>"1101100101110001",
936=>"1111101100011010",
937=>"0001000111000101",
938=>"0001000011111100",
939=>"1101100001011100",
940=>"1011101001001001",
941=>"0010111001000100",
942=>"0111111011011101",
943=>"0001110010110111",
944=>"1011110110100001",
945=>"1100100101001010",
946=>"0000010111001100",
947=>"0010011011100011",
948=>"1111110110000000",
949=>"1101100000000101",
950=>"1111001011000111",
951=>"0000111001110001",
952=>"0001010100110010",
953=>"1110101010000101",
954=>"1011010100111101",
955=>"0000101110001011",
956=>"0111110101001100",
957=>"0011110110010010",
958=>"1100101000011010",
959=>"1011111000101000",
960=>"1111011110011101",
961=>"0010011010000110",
962=>"0000101101111100",
963=>"1101101001111100",
964=>"1110100101110100",
965=>"0000101001100101",
966=>"0001011001101000",
967=>"1111101010010100",
968=>"1011100000111010",
969=>"1110101001111010",
970=>"0110111100111100",
971=>"0101100111011110",
972=>"1101111000100010",
973=>"1011100011100011",
974=>"1110011100001110",
975=>"0010000001101011",
976=>"0001100011111000",
977=>"1110000101100010",
978=>"1110000010100110",
979=>"0000010010000100",
980=>"0001010101011010",
981=>"0000011011111000",
982=>"1100010010111011",
983=>"1100111011000000",
984=>"0101011001001111",
985=>"0111000001100000",
986=>"1111011111100010",
987=>"1011011011100011",
988=>"1101100010100011",
989=>"0001011010110011",
990=>"0010001000101110",
991=>"1110110010101010",
992=>"1101101001101010",
993=>"1111110010100101",
994=>"0001001010110111",
995=>"0001000001110001",
996=>"1101010011110111",
997=>"1011110100011001",
998=>"0011011100010101",
999=>"0111110011100101",
1000=>"0001011100101100",
1001=>"1011110011011000",
1002=>"1100100110111001",
1003=>"0000011100000011",
1004=>"0010011011101001",
1005=>"1111110011100001",
1006=>"1101011100110100",
1007=>"1111001101101111",
1008=>"0000110111111101",
1009=>"0001010101111110",
1010=>"1110100011110100",
1011=>"1011010001100001",
1012=>"0000110100100111",
1013=>"0111110100000001",
1014=>"0011101110110101",
1015=>"1100100110101011",
1016=>"1011111100011110",
1017=>"1111011111011110",
1018=>"0010010111111011",
1019=>"0000101110010111",
1020=>"1101100111100100",
1021=>"1110101000101001",
1022=>"0000101001110100",
1023=>"0001011000000000");
  
  rom2 <= (
0=>"1111100101001100",
1=>"1011100010001001",
2=>"1110101111101101",
3=>"0110111110110001",
4=>"0101100001101011",
5=>"1101110011010000",
6=>"1011100010110000",
7=>"1110100010010110",
8=>"0010000010111101",
9=>"0001100010110001",
10=>"1110000101011011",
11=>"1110000100000111",
12=>"0000010100000011",
13=>"0001010101000001",
14=>"0000011000110011",
15=>"1100001111100100",
16=>"1101000000010010",
17=>"0101011111111010",
18=>"0110111110001111",
19=>"1111011001011010",
20=>"1011011101101101",
21=>"1101100110100101",
22=>"0001011101011010",
23=>"0010000111011100",
24=>"1110101111001100",
25=>"1101101001101001",
26=>"1111110011110010",
27=>"0001001001010011",
28=>"0000111111011010",
29=>"1101001101110100",
30=>"1011110111101100",
31=>"0011100001011000",
32=>"0111110101000001",
33=>"0001010010111001",
34=>"1011101011100111",
35=>"1100101111110110",
36=>"0000101001101000",
37=>"0010011001010101",
38=>"1111100111011100",
39=>"1101011101100111",
40=>"1111010101010011",
41=>"0000111011110100",
42=>"0001010000110001",
43=>"1110010110000110",
44=>"1011010011001101",
45=>"0001010110000011",
46=>"0111111010101001",
47=>"0011010011110101",
48=>"1100010110101000",
49=>"1100000111000000",
50=>"1111101100100100",
51=>"0010011011010101",
52=>"0000100010111001",
53=>"1101100101101000",
54=>"1110110001000011",
55=>"0000101100101001",
56=>"0001011000100001",
57=>"1111011001110111",
58=>"1011011011111100",
59=>"1111001100100110",
60=>"0111001111001011",
61=>"0101001010000110",
62=>"1101100001000001",
63=>"1011100111110110",
64=>"1110101111111001",
65=>"0010001001000101",
66=>"0001010101100100",
67=>"1101111101011110",
68=>"1110001010110111",
69=>"0000011001010000",
70=>"0001010111000110",
71=>"0000001111001001",
72=>"1100000000001111",
73=>"1101010110010001",
74=>"0101110111111101",
75=>"0110101100111011",
76=>"1111000100110001",
77=>"1011011001100101",
78=>"1101110110000011",
79=>"0001100011011101",
80=>"0001111111110010",
81=>"1110100011011010",
82=>"1101110000001100",
83=>"1111111001101111",
84=>"0001001011010001",
85=>"0000111100110011",
86=>"1101001011111001",
87=>"1011111011100101",
88=>"0011101010000001",
89=>"0111110011110100",
90=>"0001001100011110",
91=>"1011101001000110",
92=>"1100110010000100",
93=>"0000101110011010",
94=>"0010011010001110",
95=>"1111100010000011",
96=>"1101100000001110",
97=>"1111010110111001",
98=>"0001000000100010",
99=>"0001010010001100",
100=>"1110010001001110",
101=>"1011010100010010",
102=>"0001011110110101",
103=>"0111111011011011",
104=>"0011001001111000",
105=>"1100010101110111",
106=>"1100000111110111",
107=>"1111101110010011",
108=>"0010011110101100",
109=>"0000011101000111",
110=>"1101100011001110",
111=>"1110110000100011",
112=>"0000110000101100",
113=>"0001011000001101",
114=>"1111010101011111",
115=>"1011011010110011",
116=>"1111010001011001",
117=>"0111010011001111",
118=>"0101000011000001",
119=>"1101011010011011",
120=>"1011100111100100",
121=>"1110110011000111",
122=>"0010001100111011",
123=>"0001010010100101",
124=>"1101111010110011",
125=>"1110001100101011",
126=>"0000011000011011",
127=>"0001010110111100",
128=>"0000010000011000",
129=>"1011111111100011",
130=>"1101011110101111",
131=>"0101111111010011",
132=>"0110100111101001",
133=>"1110111100000111",
134=>"1011011011001010",
135=>"1101110101101000",
136=>"0001101000001110",
137=>"0001111011110010",
138=>"1110100001011101",
139=>"1101110011011101",
140=>"1111111110111010",
141=>"0001001101101001",
142=>"0000110110011111",
143=>"1100111000110100",
144=>"1100000110001011",
145=>"0100000111000100",
146=>"0111101010111101",
147=>"0000110000000111",
148=>"1011100100010010",
149=>"1100111111101111",
150=>"0000110111000111",
151=>"0010011011010110",
152=>"1111010111110001",
153=>"1101100001010101",
154=>"1111011110011100",
155=>"0001000010000011",
156=>"0001001101000011",
157=>"1110000010011000",
158=>"1011011001001101",
159=>"0001111100110010",
160=>"0111111110101010",
161=>"0010101011100011",
162=>"1100001001010111",
163=>"1100001111010111",
164=>"1111111101100010",
165=>"0010011101010010",
166=>"0000010011001011",
167=>"1101100001000010",
168=>"1110111001010010",
169=>"0000110001100011",
170=>"0001010111000000",
171=>"1111000101101101",
172=>"1011010110011010",
173=>"1111101110000101",
174=>"0111100001010100",
175=>"0100101000100010",
176=>"1101000111101110",
177=>"1011110000000111",
178=>"1111000000100100",
179=>"0010001110011000",
180=>"0001000110011101",
181=>"1101110100101001",
182=>"1110010111001001",
183=>"0000011110011111",
184=>"0001010111011000",
185=>"0000000010100111",
186=>"1011110110100011",
187=>"1101110101100100",
188=>"0110010110100010",
189=>"0110010110000101",
190=>"1110110001110110",
191=>"1011011011010011",
192=>"1101111001100100",
193=>"0001101010111000",
194=>"0001111001110101",
195=>"1110100000110101",
196=>"1101110001000100",
197=>"0000000001100011",
198=>"0001001011000011",
199=>"0000110101000010",
200=>"1100110110001100",
201=>"1100001010111011",
202=>"0100001111001001",
203=>"0111100111101110",
204=>"0000101001110000",
205=>"1011100011000110",
206=>"1101000100000100",
207=>"0000111000010010",
208=>"0010010111100000",
209=>"1111010101101010",
210=>"1101100010110100",
211=>"1111100000111000",
212=>"0001000001111000",
213=>"0001001101011111",
214=>"1101111110100011",
215=>"1011011100110011",
216=>"0010000100101110",
217=>"0111111100101001",
218=>"0010100111111001",
219=>"1100000111101010",
220=>"1100010010110110",
221=>"0000000001101010",
222=>"0010011101101100",
223=>"0000001101100100",
224=>"1101100001000101",
225=>"1110111010011101",
226=>"0000110101110001",
227=>"0001010111011000",
228=>"1111000010011001",
229=>"1011010010111010",
230=>"1111110111110110",
231=>"0111100001110111",
232=>"0100100110001111",
233=>"1101000110000111",
234=>"1011101110011111",
235=>"1111000110100011",
236=>"0010001111001100",
237=>"0001000101101100",
238=>"1101101111110110",
239=>"1110011001001000",
240=>"0000011101110001",
241=>"0001010111101100",
242=>"1111111111110010",
243=>"1011101111011110",
244=>"1101111010011100",
245=>"0110011001000110",
246=>"0110001111001110",
247=>"1110011111110000",
248=>"1011011100100100",
249=>"1110000111001011",
250=>"0001110001010101",
251=>"0001110011111001",
252=>"1110010110001001",
253=>"1101111000101000",
254=>"0000001000000010",
255=>"0001010000011111",
256=>"0000101011001110",
257=>"1100101000110010",
258=>"1100011100101100",
259=>"0100101001110001",
260=>"0111011010001001",
261=>"0000001101010110",
262=>"1011100000001010",
263=>"1101001101110111",
264=>"0001000110001111",
265=>"0010010011110001",
266=>"1111001001110100",
267=>"1101100010111100",
268=>"1111101000001101",
269=>"0001000111011001",
270=>"0001000111000101",
271=>"1101101110001110",
272=>"1011100011000111",
273=>"0010100010010010",
274=>"0111111101101000",
275=>"0010001001100100",
276=>"1011111110001001",
277=>"1100011100010110",
278=>"0000010000001101",
279=>"0010011111100011",
280=>"1111111111111111",
281=>"1101011101011110",
282=>"1111000010010111",
283=>"0000110100100011",
284=>"0001010110111110",
285=>"1110110100011101",
286=>"1011010011100100",
287=>"0000010110100100",
288=>"0111101110010010",
289=>"0100001010000011",
290=>"1100110011111001",
291=>"1011110100011000",
292=>"1111010011010000",
293=>"0010010101010001",
294=>"0000111000010111",
295=>"1101101101001100",
296=>"1110011011001110",
297=>"0000100000111011",
298=>"0001010111100101",
299=>"1111111100100111",
300=>"1011101100100110",
301=>"1110000000101101",
302=>"0110011111101100",
303=>"0110001100000101",
304=>"1110010111100010",
305=>"1011011101100111",
306=>"1110001010100000",
307=>"0001110110001011",
308=>"0001110100101011",
309=>"1110010011101110",
310=>"1101111010101000",
311=>"0000001000010001",
312=>"0001010001001000",
313=>"0000101001101111",
314=>"1100100110000011",
315=>"1100011110001100",
316=>"0100110011111000",
317=>"0111010111010000",
318=>"0000000100111110",
319=>"1011011111100011",
320=>"1101010000000100",
321=>"0001000111101111",
322=>"0010010001100011",
323=>"1111000110101100",
324=>"1101100100000101",
325=>"1111101000111000",
326=>"0001000101101010",
327=>"0001000110011100",
328=>"1101101001000110",
329=>"1011100100110110",
330=>"0010101001100111",
331=>"0111111101001011",
332=>"0010000000110011",
333=>"1011111010101010",
334=>"1100100000001100",
335=>"0000010000111100",
336=>"0010011011111101",
337=>"1111111100010110",
338=>"1101100000001111",
339=>"1111000111001100",
340=>"0000111000000001",
341=>"0001010101101111",
342=>"1110110001100001",
343=>"1011010101000000",
344=>"0000011110111010",
345=>"0111110001011100",
346=>"0100000011101111",
347=>"1100101111110101",
348=>"1011110100111111",
349=>"1111010111101001",
350=>"0010011000011110",
351=>"0000110011111011",
352=>"1101101100001011",
353=>"1110100001111001",
354=>"0000100111010011",
355=>"0001011001100000",
356=>"1111110000101010",
357=>"1011100100101101",
358=>"1110011100100010",
359=>"0110110100001110",
360=>"0101110010110010",
361=>"1110000010101101",
362=>"1011100001111010",
363=>"1110010101101001",
364=>"0001111101110111",
365=>"0001101000110110",
366=>"1110001001101100",
367=>"1101111111010111",
368=>"0000001111000110",
369=>"0001010100101101",
370=>"0000100000011010",
371=>"1100011001010101",
372=>"1100110001010001",
373=>"0101001100011011",
374=>"0111001001001011",
375=>"1111101100000011",
376=>"1011011100010101",
377=>"1101011100010100",
378=>"0001010101101000",
379=>"0010001011110101",
380=>"1110111000010010",
381=>"1101100111101010",
382=>"1111101111001010",
383=>"0001001001011010",
384=>"0001000100101100",
385=>"1101011011011001",
386=>"1011101111001101",
387=>"0011001100110101",
388=>"0111110111001111",
389=>"0001101000010111",
390=>"1011110001101011",
391=>"1100101000000001",
392=>"0000011110101110",
393=>"0010011100011010",
394=>"1111101101100111",
395=>"1101100000100110",
396=>"1111001111001010",
397=>"0000111011011100",
398=>"0001010011101111",
399=>"1110100000101001",
400=>"1011010000001110",
401=>"0000111110011111",
402=>"0111110101100001",
403=>"0011110111011101",
404=>"1100101111100111",
405=>"1011110111110010",
406=>"1111011001011111",
407=>"0010010101110010",
408=>"0000110100110001",
409=>"1101101001011110",
410=>"1110100100111000",
411=>"0000100111011101",
412=>"0001011000000110",
413=>"1111101011011100",
414=>"1011100101110010",
415=>"1110100010010000",
416=>"0110110110010100",
417=>"0101101101000011",
418=>"1101111101011001",
419=>"1011100000111010",
420=>"1110011011101110",
421=>"0001111111010110",
422=>"0001100111101011",
423=>"1110001001100101",
424=>"1110000000110011",
425=>"0000010001001001",
426=>"0001010100010101",
427=>"0000011101011101",
428=>"1100010101110101",
429=>"1100110110010110",
430=>"0101010011001111",
431=>"0111000110001101",
432=>"1111100101110010",
433=>"1011011110010101",
434=>"1101100000011000",
435=>"0001011000010011",
436=>"0010001010101010",
437=>"1110110100110011",
438=>"1101100111100011",
439=>"1111110000011000",
440=>"0001000111111100",
441=>"0001000010010100",
442=>"1101010101011110",
443=>"1011110001111111",
444=>"0011010010010111",
445=>"0111111000000111",
446=>"0001100000101110",
447=>"1011101111000100",
448=>"1100101010011100",
449=>"0000100011100011",
450=>"0010011010011010",
451=>"1111101101101101",
452=>"1101011101010101",
453=>"1111010001010100",
454=>"0000111010010101",
455=>"0001010001111010",
456=>"1110011101111011",
457=>"1011010001111100",
458=>"0001000110100110",
459=>"0111111000010110",
460=>"0011100001100111",
461=>"1100011101000111",
462=>"1100000010111001",
463=>"1111100110000100",
464=>"0010011010000011",
465=>"0000101001000111",
466=>"1101100111010101",
467=>"1110101101000110",
468=>"0000101010100100",
469=>"0001011000100110",
470=>"1111100000100100",
471=>"1011011110110001",
472=>"1110111110100110",
473=>"0111000111110000",
474=>"0101010110000110",
475=>"1101101010011111",
476=>"1011100101100111",
477=>"1110101001001100",
478=>"0010000101111011",
479=>"0001011010110100",
480=>"1110000001001000",
481=>"1110000111011011",
482=>"0000010110011011",
483=>"0001010110100100",
484=>"0000010100001100",
485=>"1100000110001000",
486=>"1101001011010000",
487=>"0101101100010010",
488=>"0110110101011111",
489=>"1111010000111101",
490=>"1011011001011111",
491=>"1101101111110001",
492=>"0001011110101010",
493=>"0010000011011011",
494=>"1110101000101010",
495=>"1101101101110101",
496=>"1111111001010100",
497=>"0001001010101111",
498=>"0000111100011011",
499=>"1101000100001000",
500=>"1011111100010010",
501=>"0011110000001111",
502=>"0111101110111100",
503=>"0001000101111110",
504=>"1011101001011001",
505=>"1100110110011000",
506=>"0000101101011001",
507=>"0010011001010001",
508=>"1111100001100011",
509=>"1101011100110111",
510=>"1111010011011101",
511=>"0000111110101010",
512=>"0001010011110001",
513=>"1110011000111001",
514=>"1011010010111001",
515=>"0001001111001100",
516=>"0111111001101001",
517=>"0011010111100011",
518=>"1100011100001011",
519=>"1100000011110011",
520=>"1111100111101100",
521=>"0010011101100010",
522=>"0000100011011110",
523=>"1101100100101111",
524=>"1110101100100110",
525=>"0000101110011110",
526=>"0001011000100011",
527=>"1111011100001000",
528=>"1011011101100011",
529=>"1111000011001110",
530=>"0111001100000011",
531=>"0101001111001100",
532=>"1101100011110001",
533=>"1011100101001100",
534=>"1110101100010110",
535=>"0010001001110111",
536=>"0001010111111111",
537=>"1101111110010100",
538=>"1110001001001110",
539=>"0000010101101011",
540=>"0001010110010011",
541=>"0000010101100001",
542=>"1100000101010101",
543=>"1101010011100010",
544=>"0101110011110110",
545=>"0110110000100100",
546=>"1111001000000011",
547=>"1011011011000010",
548=>"1101101111010011",
549=>"0001100011011100",
550=>"0001111111101001",
551=>"1110100110011111",
552=>"1101110001000001",
553=>"1111111011100111",
554=>"0001001100100010",
555=>"0000111001110100",
556=>"1101000000011000",
557=>"1011111111000101",
558=>"0011111000100111",
559=>"0111101111010110",
560=>"0000111101110110",
561=>"1011100110101111",
562=>"1100111010001110",
563=>"0000110001000101",
564=>"0010011101000011",
565=>"1111011101111110",
566=>"1101100000100001",
567=>"1111011010100101",
568=>"0001000000100111",
569=>"0001001110101100",
570=>"1110001010010000",
571=>"1011010110110000",
572=>"0001101101001100",
573=>"0111111101111101",
574=>"0010111001100010",
575=>"1100001110110100",
576=>"1100001011000011",
577=>"1111110110111001",
578=>"0010011100110010",
579=>"0000011001010110",
580=>"1101100010010111",
581=>"1110110101000111",
582=>"0000101111101111",
583=>"0001010111010001",
584=>"1111001100111010",
585=>"1011011000000100",
586=>"1111011111101011",
587=>"0111011010111111",
588=>"0100110101100010",
589=>"1101010000000100",
590=>"1011101101100000",
591=>"1110111001101100",
592=>"0010001011111110",
593=>"0001001011110010",
594=>"1101111000000000",
595=>"1110010011001100",
596=>"0000011100010010",
597=>"0001010110100100",
598=>"0000001000100000",
599=>"1011111011010000",
600=>"1101101010001001",
601=>"0110001011010010",
602=>"0110100000010011",
603=>"1110101111001011",
604=>"1011011001101011",
605=>"1101111101001011",
606=>"0001101111101100",
607=>"0001110111011100",
608=>"1110011101010101",
609=>"1101110100011011",
610=>"0000000011011000",
611=>"0001010000001100",
612=>"0000110011110000",
613=>"1100110001010110",
614=>"1100010000010011",
615=>"0100010101000110",
616=>"0111101010111111",
617=>"0000111000010100",
618=>"1011100100101110",
619=>"1100111111000000",
620=>"0000110010000001",
621=>"0010011001100101",
622=>"1111011011011111",
623=>"1101100010001010",
624=>"1111011100110110",
625=>"0001000000101001",
626=>"0001001110111110",
627=>"1110000110101000",
628=>"1011011001111000",
629=>"0001110101011100",
630=>"0111111100000000",
631=>"0010110101111100",
632=>"1100001100111011",
633=>"1100001110100001",
634=>"1111111010111101",
635=>"0010011101011101",
636=>"0000010011101011",
637=>"1101100010010100",
638=>"1110110110001111",
639=>"0000110011111011",
640=>"0001010111110010",
641=>"1111001001101011",
642=>"1011010100010111",
643=>"1111101001001111",
644=>"0111011011111111",
645=>"0100110010111111",
646=>"1101001110101100",
647=>"1011101011100100",
648=>"1110111111110011",
649=>"0010001100110001",
650=>"0001001011001111",
651=>"1101110011000001",
652=>"1110010101001101",
653=>"0000011011100001",
654=>"0001010110111110",
655=>"0000000101101101",
656=>"1011110100010011",
657=>"1101101110011101",
658=>"0110001110100000",
659=>"0110011001010010",
660=>"1110101010111011",
661=>"1011011011111001",
662=>"1110000000100101",
663=>"0001101101001001",
664=>"0001110111111100",
665=>"1110011011000111",
666=>"1101110101100111",
667=>"0000000101000011",
668=>"0001001111011010",
669=>"0000101111001101",
670=>"1100101111101100",
671=>"1100010100101001",
672=>"0100011011110101",
673=>"0111100000000110",
674=>"0000011010011101",
675=>"1011100010000010",
676=>"1101000111111010",
677=>"0001000000101101",
678=>"0010010101111001",
679=>"1111001111111010",
680=>"1101100001100101",
681=>"1111100100100000",
682=>"0001000101111101",
683=>"0001001001010101",
684=>"1101110101111001",
685=>"1011011111100111",
686=>"0010010010101011",
687=>"0111111110100000",
688=>"0010010111011011",
689=>"1100000010111100",
690=>"1100010111100000",
691=>"0000001001110010",
692=>"0010011111100111",
693=>"0000000110011101",
694=>"1101011101111110",
695=>"1110111110011101",
696=>"0000110010100110",
697=>"0001010111101110",
698=>"1110111011110011",
699=>"1011010100010100",
700=>"0000000111011011",
701=>"0111101001101111",
702=>"0100010111001010",
703=>"1100111011111001",
704=>"1011110000110111",
705=>"1111001100101101",
706=>"0010010010111111",
707=>"0000111110100100",
708=>"1101101111001000",
709=>"1110011011001000",
710=>"0000100010010101",
711=>"0001010100101100",
712=>"1111111011000000",
713=>"1011101010110000",
714=>"1110001000110010",
715=>"0110100100110111",
716=>"0110000110010000",
717=>"1110010010000010",
718=>"1011011110101100",
719=>"1110001110111011",
720=>"0001110101011110",
721=>"0001110000011001",
722=>"1110010011001110",
723=>"1101111000100100",
724=>"0000000100101111",
725=>"0001010000011110",
726=>"0000101101011101",
727=>"1100101101001110",
728=>"1100010101101001",
729=>"0100100110001011",
730=>"0111011101011100",
731=>"0000010010000110",
732=>"1011100001000111",
733=>"1101001010001110",
734=>"0001000010001000",
735=>"0010010011111010",
736=>"1111001100100111",
737=>"1101100010101111",
738=>"1111100101001001",
739=>"0001000100010100",
740=>"0001001000101000",
741=>"1101110000111011",
742=>"1011100000111011",
743=>"0010011010001100",
744=>"0111111110001100",
745=>"0010001110111000",
746=>"1011111111000001",
747=>"1100011011011100",
748=>"0000001010100010",
749=>"0010011100001110",
750=>"0000000010100011",
751=>"1101100000101111",
752=>"1111000011001001",
753=>"0000110110010010",
754=>"0001010110011100",
755=>"1110111000111110",
756=>"1011010101011001",
757=>"0000001111110111",
758=>"0111101101000000",
759=>"0100010001001000",
760=>"1100110111011111",
761=>"1011110001101000",
762=>"1111010000101101",
763=>"0010010110101111",
764=>"0000111001110000",
765=>"1101101110101100",
766=>"1110011101111100",
767=>"0000100101000011",
768=>"0001011001001101",
769=>"1111110110111100",
770=>"1011101000110000",
771=>"1110001111100010",
772=>"0110101010111101",
773=>"0101111101110101",
774=>"1110001101000110",
775=>"1011100000100110",
776=>"1110001111000000",
777=>"0001111001111101",
778=>"0001101101100010",
779=>"1110001110000111",
780=>"1101111100001010",
781=>"0000001100001000",
782=>"0001010011110101",
783=>"0000100100110110",
784=>"1100011111110111",
785=>"1100101000000100",
786=>"0100111111001100",
787=>"0111010000011101",
788=>"1111111000101100",
789=>"1011011101011111",
790=>"1101010110000101",
791=>"0001010000011000",
792=>"0010001110101010",
793=>"1110111110000100",
794=>"1101100101110010",
795=>"1111101011101011",
796=>"0001000111111101",
797=>"0001000111010110",
798=>"1101100011000111",
799=>"1011101010010011",
800=>"0010111101100011",
801=>"0111111001101000",
802=>"0001110110000100",
803=>"1011110101110010",
804=>"1100100010101100",
805=>"0000011000100111",
806=>"0010011100111110",
807=>"1111110100001001",
808=>"1101100000001111",
809=>"1111001011100100",
810=>"0000111001011000",
811=>"0001010101001110",
812=>"1110100111110010",
813=>"1011010000011110",
814=>"0000101101111100",
815=>"0111110100011011",
816=>"0011110110000000",
817=>"1100100111011010",
818=>"1011111100001000",
819=>"1111011100000001",
820=>"0010011011011011",
821=>"0000110010011000",
822=>"1101101001001101",
823=>"1110100110010000",
824=>"0000101000000100",
825=>"0001011000000100",
826=>"1111101001010111",
827=>"1011100011010011",
828=>"1110100110001100",
829=>"0110101111001110",
830=>"0101110111100100",
831=>"1110001000000101",
832=>"1011011111001001",
833=>"1110010101001110",
834=>"0001111011011110",
835=>"0001101100011110",
836=>"1110001101111010",
837=>"1101111101100110",
838=>"0000001110001001",
839=>"0001010011100111",
840=>"0000100001111000",
841=>"1100011100010101",
842=>"1100101100110110",
843=>"0101000110001101",
844=>"0111001101101100",
845=>"1111110010010111",
846=>"1011011111001110",
847=>"1101011010010000",
848=>"0001010011000010",
849=>"0010001101101011",
850=>"1110111010100000",
851=>"1101100101101001",
852=>"1111101100111001",
853=>"0001000110100100",
854=>"0001000100111111",
855=>"1101011101001110",
856=>"1011101100110001",
857=>"0011000011001110",
858=>"0111111010101000",
859=>"0001101110101000",
860=>"1011110010110101",
861=>"1100100101001011",
862=>"0000011101010110",
863=>"0010011011010010",
864=>"1111110011111100",
865=>"1101011101010011",
866=>"1111001101010001",
867=>"0000111000110101",
868=>"0001010010110110",
869=>"1110100101101101",
870=>"1011010001001000",
871=>"0000110111001110",
872=>"0111110101011101",
873=>"0011101111010010",
874=>"1100100011111011",
875=>"1011111110111110",
876=>"1111011111100000",
877=>"0010011000100100",
878=>"0000101111001110",
879=>"1101101001010010",
880=>"1110101001001000",
881=>"0000101000011110",
882=>"0001011000100001",
883=>"1111100111001010",
884=>"1011100001111100",
885=>"1110110000111100",
886=>"0110111111110000",
887=>"0101100001110110",
888=>"1101110100001111",
889=>"1011100011101000",
890=>"1110100010011111",
891=>"0010000010100110",
892=>"0001011111110111",
893=>"1110000101000011",
894=>"1110000100000010",
895=>"0000010011100100",
896=>"0001010101111011",
897=>"0000011001000111",
898=>"1100001100001101",
899=>"1101000000101111",
900=>"0101100000001010",
901=>"0110111101101100",
902=>"1111011101010001",
903=>"1011011001110100",
904=>"1101101001011011",
905=>"0001011001110101",
906=>"0010000110101111",
907=>"1110101110001011",
908=>"1101101011011011",
909=>"1111110110000110",
910=>"0001001001011001",
911=>"0000111111100100",
912=>"1101001011110000",
913=>"1011110110000000",
914=>"0011100001011101",
915=>"0111110010100100",
916=>"0001010011101100",
917=>"1011101100011110",
918=>"1100110000111111",
919=>"0000100111010010",
920=>"0010011010101100",
921=>"1111100111011001",
922=>"1101011110101011",
923=>"1111010101111100",
924=>"0000111110011011",
925=>"0001010000110111",
926=>"1110010100011010",
927=>"1011010110011010",
928=>"0001010100111100",
929=>"0111111001000111",
930=>"0011010000101101",
931=>"1100010111110100",
932=>"1100000101001110",
933=>"1111101110000100",
934=>"0010011100100111",
935=>"0000100100000100",
936=>"1101100111001001",
937=>"1110101000001100",
938=>"0000101100100101",
939=>"0001011000011111",
940=>"1111100010110110",
941=>"1011100000011111",
942=>"1110110101011111",
943=>"0111000100001100",
944=>"0101011011010000",
945=>"1101101101010001",
946=>"1011100011001010",
947=>"1110100101011111",
948=>"0010000110101100",
949=>"0001011101001000",
950=>"1110000010001001",
951=>"1110000101110000",
952=>"0000010010111101",
953=>"0001010101011111",
954=>"0000011010100100",
955=>"1100001011010001",
956=>"1101001000110101",
957=>"0101100111111001",
958=>"0110111001001000",
959=>"1111010100001001",
960=>"1011011011010000",
961=>"1101101000111011",
962=>"0001011110100110",
963=>"0010000011001101",
964=>"1110101011110001",
965=>"1101101110101001",
966=>"1111111000010110",
967=>"0001001011010100",
968=>"0000111101000010",
969=>"1101000111111101",
970=>"1011111000100011",
971=>"0011101001110111",
972=>"0111110011010001",
973=>"0001001011100111",
974=>"1011101001100101",
975=>"1100110100110000",
976=>"0000101011000010",
977=>"0010011110011011",
978=>"1111100100010100",
979=>"1101011111110101",
980=>"1111010110101111",
981=>"0000111111000011",
982=>"0001010000001111",
983=>"1110010010000000",
984=>"1011010100111001",
985=>"0001011101100001",
986=>"0111111100110000",
987=>"0011000111011000",
988=>"1100010100101110",
989=>"1100000110110011",
990=>"1111110000010011",
991=>"0010011011111100",
992=>"0000011111100101",
993=>"1101100011110011",
994=>"1110110001000110",
995=>"0000101101101110",
996=>"0001010111100100",
997=>"1111010011110100",
998=>"1011011010010001",
999=>"1111010001010111",
1000=>"0111010100010001",
1001=>"0101000010001000",
1002=>"1101011000111010",
1003=>"1011101010111101",
1004=>"1110110011000000",
1005=>"0010001001001011",
1006=>"0001010001001011",
1007=>"1101111011010101",
1008=>"1110001111100100",
1009=>"0000011001110000",
1010=>"0001010110000000",
1011=>"0000001101110111",
1012=>"1100000000101001",
1013=>"1101011110101010",
1014=>"0110000000000110",
1015=>"0110101001110000",
1016=>"1110111010111001",
1017=>"1011011001010011",
1018=>"1101110110101000",
1019=>"0001101011001010",
1020=>"0001111011100000",
1021=>"1110100010001101",
1022=>"1101110001111100",
1023=>"1111111111111100");
  
  rom3 <= (
0=>"0001001111010111",
1=>"0000110110111111",
2=>"1100111001010010",
3=>"1100000111101011",
4=>"0100001001100101",
5=>"0111101000100101",
6=>"0000101110010001",
7=>"1011100111000010",
8=>"1100111110001110",
9=>"0000110110011100",
10=>"0010011001011110",
11=>"1111010110000001",
12=>"1101100000001011",
13=>"1111011110000010",
14=>"0001000100001110",
15=>"0001001101000111",
16=>"1110000001110011",
17=>"1011011011100110",
18=>"0001101001001101",
19=>"0111111001101110",
20=>"0011000100100100",
21=>"1100010010001001",
22=>"1100001010100111",
23=>"1111110100000001",
24=>"0010011101001001",
25=>"0000011001101000",
26=>"1101100011110111",
27=>"1110110001111110",
28=>"0000110010000101",
29=>"0001011000000011",
30=>"1111010000110101",
31=>"1011010110001101",
32=>"1111011010110110",
33=>"0111010101100011",
34=>"0100111111100001",
35=>"1101010111100101",
36=>"1011101000110111",
37=>"1110111001000011",
38=>"0010001010000111",
39=>"0001010000101011",
40=>"1101110110011000",
41=>"1110010001011000",
42=>"0000011001001100",
43=>"0001010110001110",
44=>"0000001011011010",
45=>"1011111001011100",
46=>"1101100010110100",
47=>"0110000011100000",
48=>"0110100010111101",
49=>"1110110110010111",
50=>"1011011011011101",
51=>"1101111010000011",
52=>"0001101000110001",
53=>"0001111011110100",
54=>"1110100000001110",
55=>"1101110010110001",
56=>"0000000001111101",
57=>"0001001110010011",
58=>"0000110010111111",
59=>"1100110110110001",
60=>"1100001101000010",
61=>"0100001101101011",
62=>"0111100101011111",
63=>"0000100111101110",
64=>"1011100100001100",
65=>"1101000010000100",
66=>"0000111011000010",
67=>"0010010111110011",
68=>"1111010110000110",
69=>"1101100000011010",
70=>"1111100000101110",
71=>"0001000100100000",
72=>"0001001011011010",
73=>"1101111101100100",
74=>"1011011100100101",
75=>"0010000011000011",
76=>"0111111110110000",
77=>"0010100101010101",
78=>"1100000111111111",
79=>"1100010010110111",
80=>"0000000011010010",
81=>"0010011111011100",
82=>"0000001100111001",
83=>"1101011110101101",
84=>"1110111010100001",
85=>"0000110000101010",
86=>"0001011000010000",
87=>"1111000011000101",
88=>"1011010101011100",
89=>"1111111000100010",
90=>"0111100100100001",
91=>"0100100100001010",
92=>"1101000100001010",
93=>"1011101101101100",
94=>"1111000101111100",
95=>"0010010000110001",
96=>"0001000100010001",
97=>"1101110010000000",
98=>"1110010111010001",
99=>"0000100000000000",
100=>"0001010100010100",
101=>"0000000000110010",
102=>"1011101111100001",
103=>"1101111100001001",
104=>"0110011011000000",
105=>"0110010000100001",
106=>"1110011101010000",
107=>"1011011101010100",
108=>"1110001000101110",
109=>"0001110001000000",
110=>"0001110101001011",
111=>"1110010111001100",
112=>"1101111010001011",
113=>"0000000110110001",
114=>"0001010000001100",
115=>"0000101101000110",
116=>"1100101001010111",
117=>"1100011100111110",
118=>"0100101011011101",
119=>"0111011010000111",
120=>"0000001110001111",
121=>"1011100001000100",
122=>"1101001110010101",
123=>"0001000110000011",
124=>"0010010010001111",
125=>"1111010000101110",
126=>"1101100010010011",
127=>"1111100000111110",
128=>"0001000011001011",
129=>"0001001010100000",
130=>"1101111000110111",
131=>"1011011101011010",
132=>"0010001010110010",
133=>"0111111110100011",
134=>"0010011101000001",
135=>"1100000011101011",
136=>"1100010110111001",
137=>"0000000100000001",
138=>"0010011100010001",
139=>"0000001000110010",
140=>"1101100001011100",
141=>"1110111111000110",
142=>"0000110100100001",
143=>"0001010111000001",
144=>"1111000000010101",
145=>"1011010110001111",
146=>"0000000000111111",
147=>"0111100111111111",
148=>"0100011110010101",
149=>"1100111111100000",
150=>"1011101110011110",
151=>"1111001001110000",
152=>"0010010100110001",
153=>"0000111111011111",
154=>"1101110001011011",
155=>"1110011010000011",
156=>"0000100010101101",
157=>"0001011000110101",
158=>"1111111101000010",
159=>"1011101101001011",
160=>"1110000010111000",
161=>"0110100001001011",
162=>"0110001000100100",
163=>"1110010111110010",
164=>"1011011111100000",
165=>"1110001000011101",
166=>"0001110101110110",
167=>"0001110010000110",
168=>"1110010010101101",
169=>"1101111001000101",
170=>"0000001001000101",
171=>"0001010010111101",
172=>"0000101001000011",
173=>"1100100110100110",
174=>"1100011111010011",
175=>"0100110001101010",
176=>"0111010111001101",
177=>"0000000101100100",
178=>"1011011110111000",
179=>"1101010000000000",
180=>"0001001010111100",
181=>"0010010001010100",
182=>"1111000011111100",
183=>"1101100100001001",
184=>"1111101000000110",
185=>"0001000110100000",
186=>"0001001001110001",
187=>"1101101010111011",
188=>"1011100101110110",
189=>"0010101110001101",
190=>"0111111011011000",
191=>"0010000011111001",
192=>"1011111010000111",
193=>"1100011101100111",
194=>"0000010010010100",
195=>"0010011101011101",
196=>"1111111010100001",
197=>"1101100000010100",
198=>"1111000111101110",
199=>"0000110111100100",
200=>"0001010110001101",
201=>"1110101111010100",
202=>"1011010000011111",
203=>"0000011110100101",
204=>"0111110000101110",
205=>"0100000011011010",
206=>"1100101110110101",
207=>"1011111000011010",
208=>"1111010101011011",
209=>"0010011001011110",
210=>"0000111000100110",
211=>"1101101011010111",
212=>"1110100010011011",
213=>"0000100101110000",
214=>"0001010111111111",
215=>"1111101111101100",
216=>"1011100110110110",
217=>"1110011010011001",
218=>"0110110101111001",
219=>"0101110000111000",
220=>"1110000001100000",
221=>"1011011111111100",
222=>"1110010111110010",
223=>"0001111011111101",
224=>"0001101001100010",
225=>"1110001011010110",
226=>"1110000000000000",
227=>"0000001101000110",
228=>"0001010011001100",
229=>"0000011110111100",
230=>"1100011001011001",
231=>"1100100101000111",
232=>"0100111000000010",
233=>"0111010101010010",
234=>"1111111110101010",
235=>"1011100000110011",
236=>"1101010011111000",
237=>"0001001101111011",
238=>"0010010000001110",
239=>"1111000000100100",
240=>"1101100011101100",
241=>"1111101001100100",
242=>"0001000100111110",
243=>"0001000111101010",
244=>"1101100100110111",
245=>"1011101000001011",
246=>"0010110011110101",
247=>"0111111100101011",
248=>"0001111100011110",
249=>"1011110111000010",
250=>"1100011111111011",
251=>"0000010111001011",
252=>"0010011011110011",
253=>"1111111010010100",
254=>"1101011101011010",
255=>"1111001001010000",
256=>"0000110111001110",
257=>"0001010011101111",
258=>"1110101101010101",
259=>"1011010000110111",
260=>"0000100111110110",
261=>"0111110010000010",
262=>"0011111100110010",
263=>"1100101011001010",
264=>"1011111011001010",
265=>"1111011000111110",
266=>"0010010110110100",
267=>"0000110101010011",
268=>"1101101011011010",
269=>"1110100101001111",
270=>"0000100110010010",
271=>"0001011000011010",
272=>"1111101101100011",
273=>"1011100101100001",
274=>"1110100011100000",
275=>"0110110111010011",
276=>"0101101101010000",
277=>"1101111110010100",
278=>"1011100001110110",
279=>"1110011011110101",
280=>"0001111111000011",
281=>"0001100100110010",
282=>"1110001001001000",
283=>"1110000000110000",
284=>"0000010000101000",
285=>"0001010101001111",
286=>"0000011101110100",
287=>"1100010010100010",
288=>"1100110110101000",
289=>"0101010011101010",
290=>"0111000101011011",
291=>"1111101001110100",
292=>"1011011010011010",
293=>"1101100011001010",
294=>"0001010100111001",
295=>"0010001001110011",
296=>"1110110011110110",
297=>"1101101001001101",
298=>"1111110010110010",
299=>"0001001000000001",
300=>"0001000010100000",
301=>"1101010011011110",
302=>"1011110000001110",
303=>"0011010010011110",
304=>"0111110101101011",
305=>"0001100001011011",
306=>"1011101111111100",
307=>"1100101011100111",
308=>"0000100001001111",
309=>"0010011011101001",
310=>"1111101101110000",
311=>"1101011110010011",
312=>"1111010010000010",
313=>"0000111100110100",
314=>"0001010010001101",
315=>"1110011100000011",
316=>"1011010101001101",
317=>"0001000101100001",
318=>"0111110110111000",
319=>"0011011110011011",
320=>"1100011110010000",
321=>"1100000001001110",
322=>"1111100111010011",
323=>"0010011011101101",
324=>"0000101001001000",
325=>"1101100110010100",
326=>"1110101011000000",
327=>"0000101101011101",
328=>"0001011000000010",
329=>"1111011110011000",
330=>"1011011111010001",
331=>"1110111100011011",
332=>"0111001001010111",
333=>"0101010101000100",
334=>"1101101001010010",
335=>"1011100110001101",
336=>"1110101001111110",
337=>"0010000111101011",
338=>"0001100001001101",
339=>"1110000110101111",
340=>"1110000001111100",
341=>"0000010000100000",
342=>"0001010100010110",
343=>"0000011111101001",
344=>"1100010001001111",
345=>"1100111110101111",
346=>"0101011011011001",
347=>"0111000001011011",
348=>"1111100000010100",
349=>"1011011011111001",
350=>"1101100010100001",
351=>"0001011001101101",
352=>"0010000110011100",
353=>"1110110001010001",
354=>"1101101100010101",
355=>"1111110101000111",
356=>"0001001001111100",
357=>"0001000000001010",
358=>"1101001111100010",
359=>"1011110010100110",
360=>"0011011010110101",
361=>"0111110110101111",
362=>"0001011001010111",
363=>"1011101100110110",
364=>"1100101111010011",
365=>"0000100100111111",
366=>"0010011111011111",
367=>"1111101010110000",
368=>"1101011111010010",
369=>"1111010010111100",
370=>"0000111101010111",
371=>"0001010001101100",
372=>"1110011001101000",
373=>"1011010011100110",
374=>"0001001101110100",
375=>"0111111011000001",
376=>"0011010101000110",
377=>"1100011011000001",
378=>"1100000010101001",
379=>"1111101001101111",
380=>"0010011010110100",
381=>"0000100101110101",
382=>"1101100101011010",
383=>"1110101101001000",
384=>"0000101011101000",
385=>"0001010111110011",
386=>"1111011010100011",
387=>"1011011100111011",
388=>"1111000011001111",
389=>"0111001101000001",
390=>"0101001110011100",
391=>"1101100010000110",
392=>"1011101000100010",
393=>"1110101100011010",
394=>"0010000110000110",
395=>"0001010110100000",
396=>"1101111110110100",
397=>"1110001100000011",
398=>"0000010111000110",
399=>"0001010101011001",
400=>"0000010011000000",
401=>"1100000110010100",
402=>"1101010011100011",
403=>"0101110100100001",
404=>"0110110010110000",
405=>"1111000110111000",
406=>"1011011001001011",
407=>"1101110000001001",
408=>"0001100110011101",
409=>"0001111111010111",
410=>"1110100111010001",
411=>"1101101111100000",
412=>"1111111100100101",
413=>"0001001110010011",
414=>"0000111010010101",
415=>"1101000000110110",
416=>"1100000000100000",
417=>"0011111011001100",
418=>"0111101101000110",
419=>"0000111011110111",
420=>"1011101001011111",
421=>"1100111000110100",
422=>"0000110000010100",
423=>"0010011011010011",
424=>"1111011100000100",
425=>"1101011111100001",
426=>"1111011001111010",
427=>"0001000011000000",
428=>"0001001110011110",
429=>"1110001010001010",
430=>"1011011000001010",
431=>"0001101100000010",
432=>"0111111100100001",
433=>"0010111010101101",
434=>"1100001110001101",
435=>"1100001010101011",
436=>"1111111000111000",
437=>"0010011110111100",
438=>"0000010101111110",
439=>"1101100010001011",
440=>"1110110100010000",
441=>"0000110000001001",
442=>"0001011001011001",
443=>"1111010000101100",
444=>"1011010100110100",
445=>"1111001101101100",
446=>"0111001110000000",
447=>"0101001100001100",
448=>"1101100000100000",
449=>"1011100110100101",
450=>"1110110010001000",
451=>"0010000111011100",
452=>"0001010101110100",
453=>"1101111010000110",
454=>"1110001101011111",
455=>"0000010110111000",
456=>"0001010101010100",
457=>"0000010000111111",
458=>"1011111110110011",
459=>"1101010111100111",
460=>"0101111000000010",
461=>"0110101100001111",
462=>"1111000010000000",
463=>"1011011011010111",
464=>"1101110011100000",
465=>"0001100100010011",
466=>"0001111111011100",
467=>"1110100101100001",
468=>"1101110000000010",
469=>"1111111110110101",
470=>"0001001101001000",
471=>"0000110110100110",
472=>"1100111101111101",
473=>"1100000101111100",
474=>"0011111111001110",
475=>"0111101010011001",
476=>"0000110101000110",
477=>"1011100110101100",
478=>"1100111100010100",
479=>"0000110101010001",
480=>"0010011001011110",
481=>"1111011100010111",
482=>"1101011111011011",
483=>"1111011100111010",
484=>"0001000010111110",
485=>"0001001101010101",
486=>"1110000101001101",
487=>"1011011010000100",
488=>"0001110011011000",
489=>"0111111110011011",
490=>"0010110011001101",
491=>"1100001101011011",
492=>"1100001110010100",
493=>"1111111100110001",
494=>"0010011111000000",
495=>"0000010011010100",
496=>"1101011111101011",
497=>"1110110110100100",
498=>"0000101110101000",
499=>"0001011000101110",
500=>"1111001010001110",
501=>"1011010111000000",
502=>"1111101001110101",
503=>"0111011110110001",
504=>"0100110000111100",
505=>"1101001100101111",
506=>"1011101010101110",
507=>"1110111111001101",
508=>"0010001110010010",
509=>"0001001001111001",
510=>"1101110101000100",
511=>"1110010011011110",
512=>"0000011101100110",
513=>"0001010011110111",
514=>"0000000110011001",
515=>"1011110100100101",
516=>"1101101111111001",
517=>"0110010000101001",
518=>"0110011010011011",
519=>"1110101000101100",
520=>"1011011100010011",
521=>"1110000010011011",
522=>"0001101100100101",
523=>"0001111001011010",
524=>"1110011011111100",
525=>"1101110111011010",
526=>"0000000011101000",
527=>"0001001111010000",
528=>"0000110000110111",
529=>"1100110000100011",
530=>"1100010100101001",
531=>"0100011101110001",
532=>"0111011111110111",
533=>"0000011011100010",
534=>"1011100010110000",
535=>"1101001000100101",
536=>"0001000000011011",
537=>"0010010100000110",
538=>"1111001101101111",
539=>"1101100010100001",
540=>"1111100011001100",
541=>"0001000111000001",
542=>"0001001001101101",
543=>"1101110100010110",
544=>"1011011101000001",
545=>"0010010101011001",
546=>"0111111011011111",
547=>"0010011100100000",
548=>"1011111111110110",
549=>"1100011001000000",
550=>"0000000111010110",
551=>"0010011010101111",
552=>"0000001111110101",
553=>"1101100001101111",
554=>"1110111011100010",
555=>"0000110010010001",
556=>"0001010111110110",
557=>"1111000111001111",
558=>"1011010111110011",
559=>"1111110010000001",
560=>"0111100010101010",
561=>"0100101011001000",
562=>"1101001000000010",
563=>"1011101011010100",
564=>"1111000011000000",
565=>"0010010010011001",
566=>"0001000101010010",
567=>"1101110100001110",
568=>"1110010110010111",
569=>"0000100000001010",
570=>"0001011000100001",
571=>"0000000010110010",
572=>"1011110010000010",
573=>"1101110110011011",
574=>"0110010111000100",
575=>"0110010010110001",
576=>"1110100010111000",
577=>"1011011110100010",
578=>"1110000010000100",
579=>"0001110001011100",
580=>"0001110110100011",
581=>"1110010111010110",
582=>"1101110110010000",
583=>"0000000101110110",
584=>"0001010010000110",
585=>"0000101100111110",
586=>"1100101101100111",
587=>"1100010110111000",
588=>"0100100011111100",
589=>"0111011101010110",
590=>"0000010010101101",
591=>"1011100000011110",
592=>"1101001010000110",
593=>"0001000101010011",
594=>"0010010011110101",
595=>"1111001001110010",
596=>"1101100010110011",
597=>"1111100100010110",
598=>"0001000101001000",
599=>"0001001011111001",
600=>"1101110010110111",
601=>"1011100001110010",
602=>"0010011110111001",
603=>"0111111100011011",
604=>"0010010001110111",
605=>"1011111110101011",
606=>"1100011000110011",
607=>"0000001011110100",
608=>"0010011101110010",
609=>"0000000000110010",
610=>"1101100000101110",
611=>"1111000011101110",
612=>"0000110101110101",
613=>"0001010110111011",
614=>"1110110110111001",
615=>"1011010000110100",
616=>"0000001111011111",
617=>"0111101100010011",
618=>"0100010000110100",
619=>"1100110110011100",
620=>"1011110101000001",
621=>"1111001110101010",
622=>"0010010111011110",
623=>"0000111110100011",
624=>"1101101101111011",
625=>"1110011110011110",
626=>"0000100011100010",
627=>"0001010111101100",
628=>"1111110101111000",
629=>"1011101010111011",
630=>"1110001101011101",
631=>"0110101100100000",
632=>"0101111100000110",
633=>"1110001011110010",
634=>"1011011110101100",
635=>"1110010000111111",
636=>"0001111000010100",
637=>"0001101101111001",
638=>"1110010000000101",
639=>"1101111100011111",
640=>"0000001010100111",
641=>"0001010001101100",
642=>"0000100100010011",
643=>"1100011110001000",
644=>"1100101000011100",
645=>"0100111111011010",
646=>"0111010001001001",
647=>"1111110110000111",
648=>"1011011111100110",
649=>"1101011000001100",
650=>"0001001101000011",
651=>"0010001100010010",
652=>"1110111101110001",
653=>"1101101000001101",
654=>"1111101101101010",
655=>"0001001000010101",
656=>"0001000011111110",
657=>"1101100101110111",
658=>"1011100100111101",
659=>"0010100011111011",
660=>"0111111110011000",
661=>"0010001010001101",
662=>"1011111011101011",
663=>"1100011010110000",
664=>"0000010000111100",
665=>"0010011100000110",
666=>"0000000000101011",
667=>"1101011101101110",
668=>"1111000101001111",
669=>"0000110101100011",
670=>"0001010100011110",
671=>"1110110100111001",
672=>"1011010001000011",
673=>"0000011000100111",
674=>"0111101110000001",
675=>"0100001010001011",
676=>"1100110010101011",
677=>"1011110111100011",
678=>"1111010010011010",
679=>"0010010100110101",
680=>"0000111011010010",
681=>"1101101101110010",
682=>"1110100001010111",
683=>"0000100100000011",
684=>"0001011000001010",
685=>"1111110011110011",
686=>"1011101001011100",
687=>"1110010110011001",
688=>"0110101110010100",
689=>"0101111000010110",
690=>"1110001000101011",
691=>"1011100000010011",
692=>"1110010101001110",
693=>"0001111011010100",
694=>"0001101001100010",
695=>"1110001101011010",
696=>"1101111101100101",
697=>"0000001101100111",
698=>"0001010100011101",
699=>"0000100010010100",
700=>"1100011001000110",
701=>"1100101100111011",
702=>"0101000110110011",
703=>"0111001100101101",
704=>"1111110110100010",
705=>"1011011011010011",
706=>"1101011100111101",
707=>"0001001111110010",
708=>"0010001100101010",
709=>"1110111001101000",
710=>"1101100111001000",
711=>"1111101111011010",
712=>"0001000110101001",
713=>"0001000101001111",
714=>"1101011011010000",
715=>"1011101010111011",
716=>"0011000011010111",
717=>"0111111000001100",
718=>"0001101111010000",
719=>"1011110011101111",
720=>"1100100110010111",
721=>"0000011011000110",
722=>"0010011100011001",
723=>"1111110100000111",
724=>"1101011110001011",
725=>"1111001110000011",
726=>"0000111011001101",
727=>"0001010011011000",
728=>"1110100011101011",
729=>"1011010100011011",
730=>"0000110110001100",
731=>"0111110100000010",
732=>"0011101100000011",
733=>"1100100101000001",
734=>"1011111101011001",
735=>"1111100000100101",
736=>"0010011010010101",
737=>"0000101111001101",
738=>"1101101000011000",
739=>"1110100110111011",
740=>"0000101011010100",
741=>"0001011000000111",
742=>"1111100100111010",
743=>"1011100010011100",
744=>"1110101110110010",
745=>"0111000001001111",
746=>"0101100001000001",
747=>"1101110010110011",
748=>"1011100100011101",
749=>"1110100010111001",
750=>"0010000100111111",
751=>"0001100000001000",
752=>"1110000010101011",
753=>"1110000011101111",
754=>"0000010000010000",
755=>"0001010011100010",
756=>"0000011011010001",
757=>"1100001101000001",
758=>"1101000011001111",
759=>"0101100000111000",
760=>"0110111111010101",
761=>"1111011000100011",
762=>"1011011011010001",
763=>"1101100100111111",
764=>"0001010100111010",
765=>"0010001001100001",
766=>"1110110110110100",
767=>"1101101010010001",
768=>"1111110001101101",
769=>"0001001000101001",
770=>"0001000010111111",
771=>"1101010111010010",
772=>"1011101101000010",
773=>"0011001011110001",
774=>"0111111001100001",
775=>"0001100111010100",
776=>"1011110000010101",
777=>"1100101010000011",
778=>"0000011110110001",
779=>"0010100000011000",
780=>"1111110001001011",
781=>"1101011111000001",
782=>"1111001111000010",
783=>"0000111011101110",
784=>"0001010010111011",
785=>"1110100001010001",
786=>"1011010010101100",
787=>"0000111110010001",
788=>"0111111000100110",
789=>"0011100010110100",
790=>"1100100001100100",
791=>"1011111110101111",
792=>"1111100011000011",
793=>"0010011001100010",
794=>"0000101011111100",
795=>"1101100111010100",
796=>"1110101001000111",
797=>"0000101001100001",
798=>"0001010111110110",
799=>"1111100001001100",
800=>"1011011111111000",
801=>"1110110101011100",
802=>"0111000101001011",
803=>"0101011010100011",
804=>"1101101011100011",
805=>"1011100110011010",
806=>"1110100101110000",
807=>"0010000010111001",
808=>"0001011011100111",
809=>"1110000010100011",
810=>"1110001000100100",
811=>"0000010100011100",
812=>"0001010100101010",
813=>"0000011000000010",
814=>"1100001100001010",
815=>"1101001000111011",
816=>"0101101000011110",
817=>"0110111011011001",
818=>"1111010011000000",
819=>"1011011001011010",
820=>"1101101001101001",
821=>"0001100001101100",
822=>"0010000010111100",
823=>"1110101100100011",
824=>"1101101101001010",
825=>"1111111001001110",
826=>"0001001101000111",
827=>"0000111101100100",
828=>"1101001000011001",
829=>"1011111001111100",
830=>"0011101100011101",
831=>"0111110001001100",
832=>"0001001001011100",
833=>"1011101100010111",
834=>"1100110011011001",
835=>"0000101010010000",
836=>"0010011100101101",
837=>"1111100010011001",
838=>"1101011110110011",
839=>"1111010110000100",
840=>"0001000001010110",
841=>"0001010000001101",
842=>"1110010001101101",
843=>"1011010110011111",
844=>"0001011100001110",
845=>"0111111011100100",
846=>"0011000111111100",
847=>"1100010110101110",
848=>"1100000111101000",
849=>"1111110001101011",
850=>"0010011110100100",
851=>"0000011100000000",
852=>"1101100011101111",
853=>"1110110000000111",
854=>"0000101110001011",
855=>"0001011001100111",
856=>"1111010111011100",
857=>"1011011001110101",
858=>"1111010110010011",
859=>"0111010100000001",
860=>"0101000011000111",
861=>"1101011010111101",
862=>"1011100111110100",
863=>"1110110011000011",
864=>"0010001011010110",
865=>"0001010000010001",
866=>"1101111010010010",
867=>"1110010000011100",
868=>"0000011001011111",
869=>"0001010101110110",
870=>"0000001111010000",
871=>"1100000111101110",
872=>"1101001101000010",
873=>"0101101100000110",
874=>"0110110101001011",
875=>"1111001101101101",
876=>"1011011110011101",
877=>"1101101101100010",
878=>"0001011111011000",
879=>"0010000011000110",
880=>"1110101010110001",
881=>"1101101101100111",
882=>"1111111011011111",
883=>"0001001100000011",
884=>"0000111001110110",
885=>"1101000101011010",
886=>"1011111111001011",
887=>"0011110000101100",
888=>"0111101110100111",
889=>"0001000010101101",
890=>"1011101001011001",
891=>"1100110110110000",
892=>"0000101111010100",
893=>"0010011010111111",
894=>"1111100010100100",
895=>"1101011110110001",
896=>"1111011000111100",
897=>"0001000001100000",
898=>"0001001111000000",
899=>"1110001100111011",
900=>"1011010111111100",
901=>"0001100011110100",
902=>"0111111101011001",
903=>"0011000001001000",
904=>"1100010011000101",
905=>"1100001010000010",
906=>"1111110110000110",
907=>"0010011110011100",
908=>"0000011001100111",
909=>"1101100000111101",
910=>"1110110010100010",
911=>"0000101100101011",
912=>"0001011000111011",
913=>"1111010001010101",
914=>"1011011000111010",
915=>"1111011011011010",
916=>"0111011000010110",
917=>"0100111101100111",
918=>"1101010101100010",
919=>"1011101000000011",
920=>"1110111000010110",
921=>"0010001011101110",
922=>"0001001111010001",
923=>"1101111000011101",
924=>"1110001111101001",
925=>"0000011011001111",
926=>"0001010011001110",
927=>"0000001011111010",
928=>"1011111001110110",
929=>"1101100100000111",
930=>"0110000101101110",
931=>"0110100100000101",
932=>"1110110100010000",
933=>"1011011011101100",
934=>"1101111100000010",
935=>"0001101000001001",
936=>"0001111101010100",
937=>"1110100000111111",
938=>"1101110100101000",
939=>"0000000000100100",
940=>"0001001110000111",
941=>"0000110100100100",
942=>"1100110111101110",
943=>"1100001100111110",
944=>"0100001111101000",
945=>"0111100101010001",
946=>"0000101000110001",
947=>"1011100100111011",
948=>"1101000010110000",
949=>"0000111010110001",
950=>"0010010110000101",
951=>"1111010011110100",
952=>"1101100001010111",
953=>"1111011111011011",
954=>"0001000101100000",
955=>"0001001011110100",
956=>"1101111100000110",
957=>"1011011001111001",
958=>"0010000101110000",
959=>"0111111011110101",
960=>"0010101010001001",
961=>"1100000101011010",
962=>"1100010011100111",
963=>"0000000010101101",
964=>"0010011100100010",
965=>"0000001100110000",
966=>"1101011110100110",
967=>"1110111101100111",
968=>"0000110001010001",
969=>"0001011000010010",
970=>"1111000010110011",
971=>"1011010101110010",
972=>"1111111000000101",
973=>"0111100011000111",
974=>"0100100010111100",
975=>"1101000110011000",
976=>"1011110001010000",
977=>"1110111101100111",
978=>"0010001111011110",
979=>"0001001011001000",
980=>"1101110111001000",
981=>"1110010010110101",
982=>"0000011101011011",
983=>"0001011000010100",
984=>"0000000111111101",
985=>"1011111010001000",
986=>"1101101011000001",
987=>"0110001100001011",
988=>"0110011100110100",
989=>"1110101110000101",
990=>"1011011101111100",
991=>"1101111011101001",
992=>"0001101100111000",
993=>"0001111010111001",
994=>"1110011011111100",
995=>"1101110110011011",
996=>"0000000011001010",
997=>"0001010000110110",
998=>"0000110000111101",
999=>"1100110100100011",
1000=>"1100001111001000",
1001=>"0100010101110001",
1002=>"0111100011000111",
1003=>"0000011111111010",
1004=>"1011100101011011",
1005=>"1101000111000111",
1006=>"0001000000001000",
1007=>"0010010101101101",
1008=>"1111010000000110",
1009=>"1101100001010010",
1010=>"1111100000111011",
1011=>"0001000011010011",
1012=>"0001001110010010",
1013=>"1101111010010100",
1014=>"1011011110111100",
1015=>"0010001101111000",
1016=>"0111111010100111",
1017=>"0010100000010110",
1018=>"1100000011010111",
1019=>"1100010100001101",
1020=>"0000000101010000",
1021=>"0010011101110110",
1022=>"0000000111001000",
1023=>"1101100001001110");
  
  rom4 <= (
0=>"1110111111111000",
1=>"0000110011110100",
2=>"0001010111110110",
3=>"1110111101101111",
4=>"1011010100000101",
5=>"0000000001111100",
6=>"0111100110101111",
7=>"0100011110011001",
8=>"1100111110001000",
9=>"1011110010000000",
10=>"1111000111101111",
11=>"0010010101010110",
12=>"0001000100010011",
13=>"1101110000110010",
14=>"1110011010100000",
15=>"0000100001010011",
16=>"0001010111010010",
17=>"1111111011111010",
18=>"1011101111010101",
19=>"1110000000111000",
20=>"0110100010100111",
21=>"0110000110111110",
22=>"1110010110010111",
23=>"1011011101101001",
24=>"1110001010010011",
25=>"0001110100011010",
26=>"0001110010001100",
27=>"1110010100110101",
28=>"1101111001010101",
29=>"0000000111101111",
30=>"0001010000101000",
31=>"0000101000101001",
32=>"1100100100101111",
33=>"1100011111110001",
34=>"0100110001101110",
35=>"0111011000000101",
36=>"0000000010110111",
37=>"1011100000111111",
38=>"1101010010000100",
39=>"0001000111111000",
40=>"0010001110101001",
41=>"1111000011110110",
42=>"1101100110001010",
43=>"1111101010100110",
44=>"0001000110010001",
45=>"0001000111100110",
46=>"1101101010001011",
47=>"1011100111010101",
48=>"0010101100110001",
49=>"0111111000100111",
50=>"0010000011100101",
51=>"1011111000010100",
52=>"1100011100111000",
53=>"0000010101100010",
54=>"0010011110000010",
55=>"1111111010111100",
56=>"1101011111101110",
57=>"1111000111001001",
58=>"0000111001110000",
59=>"0001010111011100",
60=>"1110111011101101",
61=>"1011010010000010",
62=>"0000001001010001",
63=>"0111101001101001",
64=>"0100010111001100",
65=>"1100111010101101",
66=>"1011110011111111",
67=>"1111001011111100",
68=>"0010010010100010",
69=>"0001000001010010",
70=>"1101110000010000",
71=>"1110011101101010",
72=>"0000100001100111",
73=>"0001010111111111",
74=>"1111111001101101",
75=>"1011101101111000",
76=>"1110001001011001",
77=>"0110100101000100",
78=>"0110000010110111",
79=>"1110010011101001",
80=>"1011011110100100",
81=>"1110001111010110",
82=>"0001110101000110",
83=>"0001101100011111",
84=>"1110010010011000",
85=>"1101111010010000",
86=>"0000001010101100",
87=>"0001010011100100",
88=>"0000100110100100",
89=>"1100100010110100",
90=>"1100100100000010",
91=>"0100111001011100",
92=>"0111010011100111",
93=>"0000000011010111",
94=>"1011011100100101",
95=>"1101010110110010",
96=>"0001001010100110",
97=>"0010001111010010",
98=>"1110111111100001",
99=>"1101100101010010",
100=>"1111101011110110",
101=>"0001000101011100",
102=>"0001000111010011",
103=>"1101100100111111",
104=>"1011101000001111",
105=>"0010110011001011",
106=>"0111111010111100",
107=>"0001111100001010",
108=>"1011111010010001",
109=>"1100100010110110",
110=>"0000010100011000",
111=>"0010011101001010",
112=>"1111111010010100",
113=>"1101011110011001",
114=>"1111001001111010",
115=>"0000111001101010",
116=>"0001010100010010",
117=>"1110101011010100",
118=>"1011010100000000",
119=>"0000100111000110",
120=>"0111110000011011",
121=>"0011111001110100",
122=>"1100101011110000",
123=>"1011111010010101",
124=>"1111010111111011",
125=>"0010010110101011",
126=>"0000110101111011",
127=>"1101101010001101",
128=>"1110100011001101",
129=>"0000101000111000",
130=>"0001011000010000",
131=>"1111101011001011",
132=>"1011100101111110",
133=>"1110100001101101",
134=>"0110110110111011",
135=>"0101101010010101",
136=>"1101111101110111",
137=>"1011100001110010",
138=>"1110011101000111",
139=>"0010000000010011",
140=>"0001100111011100",
141=>"1110001000001100",
142=>"1110000010110111",
143=>"0000001110011010",
144=>"0001010010010000",
145=>"0000100000001101",
146=>"1100010011001101",
147=>"1100111001001100",
148=>"0101010100011001",
149=>"0111000111000100",
150=>"1111100101010110",
151=>"1011011011010010",
152=>"1101100000010110",
153=>"0001010111110100",
154=>"0010000111101000",
155=>"1110110110001001",
156=>"1101101010100111",
157=>"1111110100101100",
158=>"0001000110010010",
159=>"0001000001011111",
160=>"1101010100010100",
161=>"1011110000111111",
162=>"0011010100011100",
163=>"0111110111110001",
164=>"0001011111110101",
165=>"1011101111011101",
166=>"1100100101010010",
167=>"0000011000011010",
168=>"0010100000111111",
169=>"1111110111101101",
170=>"1101011110110111",
171=>"1111001011010000",
172=>"0000111001110101",
173=>"0001010100010011",
174=>"1110101000011110",
175=>"1011010010111000",
176=>"0000101100111111",
177=>"0111110011011011",
178=>"0011110001000101",
179=>"1100101000000011",
180=>"1011111011010010",
181=>"1111011100001001",
182=>"0010011000001101",
183=>"0000110001110100",
184=>"1101101001100110",
185=>"1110100101000000",
186=>"0000100111011110",
187=>"0001010111101101",
188=>"1111100111110010",
189=>"1011100011001001",
190=>"1110101000000000",
191=>"0110111100101111",
192=>"0101100110011011",
193=>"1101110101001110",
194=>"1011100100100110",
195=>"1110011111000001",
196=>"0001111111100110",
197=>"0001100000011110",
198=>"1110000110100111",
199=>"1110000101000011",
200=>"0000010001110110",
201=>"0001010011101100",
202=>"0000011101000101",
203=>"1100010001111010",
204=>"1100111111011001",
205=>"0101011001010100",
206=>"0110111110110110",
207=>"1111100001100010",
208=>"1011011100110101",
209=>"1101100101100100",
210=>"0001011100000110",
211=>"0010000110110010",
212=>"1110110001100100",
213=>"1101101011010111",
214=>"1111110101011000",
215=>"0001001100010111",
216=>"0000111111111001",
217=>"1101010001111101",
218=>"1011110110001000",
219=>"0011011010001001",
220=>"0111110100001111",
221=>"0001010111011001",
222=>"1011101111010011",
223=>"1100101110011001",
224=>"0000100011101111",
225=>"0010011110011000",
226=>"1111100111111111",
227=>"1101100000011110",
228=>"1111010011111100",
229=>"0000111111001011",
230=>"0001010001111100",
231=>"1110011001001101",
232=>"1011010101001100",
233=>"0001001100101100",
234=>"0111111001100100",
235=>"0011010101111111",
236=>"1100011100010101",
237=>"1100000101101110",
238=>"1111101100110000",
239=>"0010011100111111",
240=>"0000100010100010",
241=>"1101100101010110",
242=>"1110101111100000",
243=>"0000101011011100",
244=>"0001011010001001",
245=>"1111011101111011",
246=>"1011011100110000",
247=>"1111000111110010",
248=>"0111001010000011",
249=>"0101001111001101",
250=>"1101100100010010",
251=>"1011100101101110",
252=>"1110101111100100",
253=>"0010000111101000",
254=>"0001010110001100",
255=>"1101111101001101",
256=>"1110001101011101",
257=>"0000010110001110",
258=>"0001010110001100",
259=>"0000010001100110",
260=>"1100000101110100",
261=>"1101010101001001",
262=>"0101110001011111",
263=>"0110110000100011",
264=>"1111000111111010",
265=>"1011011100110100",
266=>"1101110001001111",
267=>"0001100001101000",
268=>"0010000011011011",
269=>"1110101000001111",
270=>"1101101111011101",
271=>"1111111011110101",
272=>"0001001100111110",
273=>"0000111100110111",
274=>"1101001100111001",
275=>"1011111000111111",
276=>"0011100001110111",
277=>"0111110010011100",
278=>"0001010000000110",
279=>"1011101101110110",
280=>"1100110100000110",
281=>"0000100101010110",
282=>"0010011100011011",
283=>"1111101000001001",
284=>"1101100000010100",
285=>"1111010110111000",
286=>"0000111111011100",
287=>"0001010000101111",
288=>"1110010100100010",
289=>"1011010110001110",
290=>"0001010100100100",
291=>"0111111000111000",
292=>"0011001110011000",
293=>"1100011001011000",
294=>"1100000101101110",
295=>"1111101111100011",
296=>"0010011101011001",
297=>"0000100010000001",
298=>"1101100110000101",
299=>"1110110010101010",
300=>"0000101010000000",
301=>"0001011001011011",
302=>"1111011000000010",
303=>"1011011011011011",
304=>"1111001101000010",
305=>"0111001110011001",
306=>"0101001001111100",
307=>"1101011110101111",
308=>"1011100101100100",
309=>"1110110001100001",
310=>"0010001000111111",
311=>"0001010100010110",
312=>"1101111100110001",
313=>"1110001110111100",
314=>"0000010111111100",
315=>"0001010011001101",
316=>"0000010000011101",
317=>"1100000010101001",
318=>"1101011001000111",
319=>"0101111010010100",
320=>"0110101101010011",
321=>"1111000000001001",
322=>"1011011011001101",
323=>"1101110101110011",
324=>"0001100011011010",
325=>"0010000001001011",
326=>"1110100110000011",
327=>"1101110010001010",
328=>"1111111101010000",
329=>"0001001101000111",
330=>"0000110111111000",
331=>"1100111111010001",
332=>"1100000101011111",
333=>"0100000001101000",
334=>"0111101001100010",
335=>"0000110011011001",
336=>"1011100111010110",
337=>"1100111101011000",
338=>"0000110100000111",
339=>"0010010101000100",
340=>"1111011010011000",
341=>"1101100000010010",
342=>"1111011011100101",
343=>"0001000100001001",
344=>"0001001101010000",
345=>"1110000110000100",
346=>"1011011100001100",
347=>"0001110101001011",
348=>"0111111100010010",
349=>"0010110110111101",
350=>"1100001101101001",
351=>"1100010000010000",
352=>"1111111011111011",
353=>"0010011100010001",
354=>"0000010010111111",
355=>"1101011111101100",
356=>"1110111001011010",
357=>"0000101111101010",
358=>"0001011000001001",
359=>"1111001100110000",
360=>"1011011000010001",
361=>"1111101001000001",
362=>"0111011101100100",
363=>"0100101111100111",
364=>"1101001110110010",
365=>"1011101110110100",
366=>"1110111101101010",
367=>"0010001101110011",
368=>"0001001011001010",
369=>"1101110100111101",
370=>"1110010100111010",
371=>"0000011110101001",
372=>"0001010110100001",
373=>"0000000011100010",
374=>"1011110110110111",
375=>"1101110000101000",
376=>"0110001111001010",
377=>"0110010111100101",
378=>"1110101000000010",
379=>"1011011100000010",
380=>"1101110101011100",
381=>"0001101000001010",
382=>"0001111110111000",
383=>"1110100011111001",
384=>"1101110100000110",
385=>"1111111111101101",
386=>"0001010000000001",
387=>"0000110100010110",
388=>"1100111100000000",
389=>"1100000111100001",
390=>"0100000111101011",
391=>"0111101000000011",
392=>"0000101101100001",
393=>"1011100111010101",
394=>"1101000001101111",
395=>"0000111001111101",
396=>"0010011000001101",
397=>"1111010101011010",
398=>"1101100010001000",
399=>"1111011111001101",
400=>"0001000001010001",
401=>"0001010000010101",
402=>"1110000010001001",
403=>"1011011011111001",
404=>"0001111110100101",
405=>"0111111010010100",
406=>"0010101110100010",
407=>"1100001000000101",
408=>"1100010001011001",
409=>"0000000000111000",
410=>"0010011100111010",
411=>"0000001101111000",
412=>"1101100001101101",
413=>"1110111100001000",
414=>"0000110001110001",
415=>"0001011000011010",
416=>"1111000101010011",
417=>"1011011000100101",
418=>"1111110010011111",
419=>"0111011110111010",
420=>"0100101010001101",
421=>"1101001001110010",
422=>"1011101111010101",
423=>"1111000001011101",
424=>"0010001110001110",
425=>"0001000111101001",
426=>"1101110100011111",
427=>"1110010110010010",
428=>"0000011111001000",
429=>"0001010110110010",
430=>"0000000001100010",
431=>"1011110110100100",
432=>"1101110101110111",
433=>"0110010010100110",
434=>"0110010000010100",
435=>"1110100001011111",
436=>"1011011100101111",
437=>"1110000011101111",
438=>"0001110000001101",
439=>"0001110110011110",
440=>"1110011001011000",
441=>"1101111001000101",
442=>"0000000101101010",
443=>"0001001111000000",
444=>"0000101101001111",
445=>"1100101011000001",
446=>"1100011000010001",
447=>"0100100000111101",
448=>"0111011101100001",
449=>"0000010000001010",
450=>"1011100010011100",
451=>"1101001100001111",
452=>"0001000010011010",
453=>"0010010000111101",
454=>"1111001001110100",
455=>"1101100100100101",
456=>"1111100111000101",
457=>"0001000100101110",
458=>"0001001010000000",
459=>"1101110001110000",
460=>"1011100011100101",
461=>"0010011101001100",
462=>"0111111010000010",
463=>"0010010001000001",
464=>"1100000010011000",
465=>"1100011100010010",
466=>"0000001110110011",
467=>"0010011110011111",
468=>"0000000001001110",
469=>"1101100000000101",
470=>"1111000011001100",
471=>"0000110111111011",
472=>"0001010111101111",
473=>"1110110111011111",
474=>"1011010101001110",
475=>"0000001111111100",
476=>"0111100111100100",
477=>"0100001101010110",
478=>"1100111000010101",
479=>"1011110101011000",
480=>"1111001101001100",
481=>"0010010110010111",
482=>"0000111100111111",
483=>"1101110000000111",
484=>"1110100000000000",
485=>"0000100011000110",
486=>"0001010111010100",
487=>"1111111111100101",
488=>"1011110010101001",
489=>"1101111100101000",
490=>"0110011011101100",
491=>"0110001011100101",
492=>"1110011100011000",
493=>"1011011110000100",
494=>"1110001000100101",
495=>"0001110001000111",
496=>"0001110000111100",
497=>"1110010110100011",
498=>"1101111010001110",
499=>"0000001000001100",
500=>"0001010010101010",
501=>"0000101010010010",
502=>"1100101011000100",
503=>"1100011101010101",
504=>"0100101000000101",
505=>"0111011011001111",
506=>"0000001111011010",
507=>"1011100001110011",
508=>"1101010000011110",
509=>"0001000101100101",
510=>"0010010001011001",
511=>"1111000101110010",
512=>"1101100011010100",
513=>"1111101000100111",
514=>"0001000011101101",
515=>"0001001001111101",
516=>"1101101111110101",
517=>"1011100011110010",
518=>"0010100100010000",
519=>"0111111001101100",
520=>"0010001000111010",
521=>"1011111111001101",
522=>"1100011101100001",
523=>"0000001110011100",
524=>"0010011101000110",
525=>"0000000000111111",
526=>"1101011110011010",
527=>"1111000110001010",
528=>"0000110111101010",
529=>"0001010101011100",
530=>"1110110010100001",
531=>"1011010100011001",
532=>"0000010111101111",
533=>"0111101100101100",
534=>"0100000110110101",
535=>"1100110011110011",
536=>"1011111001101110",
537=>"1111010001000010",
538=>"0010010100110111",
539=>"0000111011101101",
540=>"1101101101000111",
541=>"1110100010010110",
542=>"0000100110000100",
543=>"0001011000100001",
544=>"1111110001000011",
545=>"1011101010001011",
546=>"1110010100010110",
547=>"0110101110001101",
548=>"0101110101001101",
549=>"1110001000011101",
550=>"1011011111110111",
551=>"1110010111000100",
552=>"0001111010100111",
553=>"0001101001111111",
554=>"1110001110001100",
555=>"1110000010000010",
556=>"0000001011000110",
557=>"0001010001101001",
558=>"0000100100010101",
559=>"1100011100101111",
560=>"1100110000001011",
561=>"0101000101011011",
562=>"0111001011001000",
563=>"1111110000100100",
564=>"1011011111011011",
565=>"1101011010011110",
566=>"0001010010011101",
567=>"0010001010110011",
568=>"1110111011100001",
569=>"1101101000111010",
570=>"1111110000111100",
571=>"0001000101011110",
572=>"0001000011011010",
573=>"1101011110000011",
574=>"1011101101110000",
575=>"0011000100010001",
576=>"0111110101010000",
577=>"0001101100110110",
578=>"1011110100100000",
579=>"1100101010100100",
580=>"0000011010011000",
581=>"0010011101011011",
582=>"1111110101000010",
583=>"1101011111110110",
584=>"1111001110000100",
585=>"0000111001101110",
586=>"0001010100111011",
587=>"1110100100110001",
588=>"1011010100110000",
589=>"0000110111000001",
590=>"0111110101110010",
591=>"0011101000100001",
592=>"1100101000011100",
593=>"1011111000111010",
594=>"1111010100110001",
595=>"0010010110111101",
596=>"0000110111010010",
597=>"1101101100101000",
598=>"1110100011110111",
599=>"0000100101000111",
600=>"0001010111100100",
601=>"1111101110001010",
602=>"1011100110110011",
603=>"1110011010110011",
604=>"0110110000101001",
605=>"0101110010001001",
606=>"1101111111001000",
607=>"1011100011000011",
608=>"1110011000010010",
609=>"0001111100001001",
610=>"0001100101001000",
611=>"1110001010111001",
612=>"1110000001100110",
613=>"0000001111001110",
614=>"0001010010101010",
615=>"0000100001111000",
616=>"1100011000000011",
617=>"1100110101110100",
618=>"0101001100011100",
619=>"0111000110110001",
620=>"1111101101100000",
621=>"1011100000110011",
622=>"1101011111100110",
623=>"0001010110111110",
624=>"0010001001111001",
625=>"1110110111001011",
626=>"1101101001001110",
627=>"1111110010000010",
628=>"0001001010111001",
629=>"0001000010111111",
630=>"1101011001010010",
631=>"1011110001000110",
632=>"0011001010001101",
633=>"0111110100010001",
634=>"0001100101110101",
635=>"1011110010001111",
636=>"1100101010011111",
637=>"0000100000010011",
638=>"0010011101111110",
639=>"1111110001001001",
640=>"1101100001010101",
641=>"1111001111110101",
642=>"0000111101011111",
643=>"0001010011011101",
644=>"1110100000010011",
645=>"1011010110000110",
646=>"0000111111100001",
647=>"0111110011100000",
648=>"0011100011011010",
649=>"1100100010111111",
650=>"1100000001101000",
651=>"1111100110011011",
652=>"0010011000110011",
653=>"0000101000010000",
654=>"1101100111010010",
655=>"1110101011011100",
656=>"0000101001011001",
657=>"0001011010000111",
658=>"1111100100100111",
659=>"1011011111110001",
660=>"1110111001110110",
661=>"0111000010100111",
662=>"0101011010101010",
663=>"1101101110110101",
664=>"1011100110010101",
665=>"1110101000010101",
666=>"0010000100101111",
667=>"0001011011001101",
668=>"1110000000111111",
669=>"1110001001111010",
670=>"0000010011100110",
671=>"0001010101011110",
672=>"0000010110100111",
673=>"1100001011101100",
674=>"1101001010010101",
675=>"0101100101111110",
676=>"0110110100000001",
677=>"1111010010001011",
678=>"1011011101100011",
679=>"1101101010101011",
680=>"0001011100110101",
681=>"0010000011011111",
682=>"1110101110001001",
683=>"1101101100101101",
684=>"1111111000110111",
685=>"0001001011011011",
686=>"0000111011101100",
687=>"1101001010111100",
688=>"1011111111011100",
689=>"0011101000011011",
690=>"0111101101111100",
691=>"0001001000000000",
692=>"1011101010011010",
693=>"1100110011111100",
694=>"0000101010101110",
695=>"0010011011000011",
696=>"1111100100100011",
697=>"1101100000111000",
698=>"1111011000001110",
699=>"0000111101011101",
700=>"0001010010011001",
701=>"1110011011111100",
702=>"1011010101001111",
703=>"0001000100111100",
704=>"0111110110110111",
705=>"0011011011111001",
706=>"1100011111111100",
707=>"1100000001011111",
708=>"1111101001010000",
709=>"0010011001010100",
710=>"0000100111100110",
711=>"1101101000000101",
712=>"1110101110011100",
713=>"0000101000010100",
714=>"0001011000111101",
715=>"1111011111101110",
716=>"1011100000110110",
717=>"1110111111000000",
718=>"0111000101111111",
719=>"0101010000001111",
720=>"1101101001010011",
721=>"1011100101111100",
722=>"1110101010011000",
723=>"0010000110001000",
724=>"0001011001011001",
725=>"1110000000100100",
726=>"1110001011001111",
727=>"0000010101100101",
728=>"0001010010010000",
729=>"0000010101110100",
730=>"1100000111111110",
731=>"1101001110111110",
732=>"0101101100000011",
733=>"0110110001100010",
734=>"1111001100100001",
735=>"1011011101100011",
736=>"1101110000100100",
737=>"0001011110000011",
738=>"0010000101001001",
739=>"1110101011000000",
740=>"1101110000000001",
741=>"1111111001110000",
742=>"0001001100001001",
743=>"0000111010111111",
744=>"1101000110110100",
745=>"1011111110110000",
746=>"0011110010101001",
747=>"0111101010101011",
748=>"0001000001101010",
749=>"1011101100100000",
750=>"1100111000100000",
751=>"0000101101100111",
752=>"0010010111010101",
753=>"1111011111100010",
754=>"1101100001101011",
755=>"1111011001100010",
756=>"0001000010001111",
757=>"0001001111000011",
758=>"1110001101110000",
759=>"1011011010000001",
760=>"0001100011000111",
761=>"0111111001111000",
762=>"0011000010010010",
763=>"1100010011101010",
764=>"1100001011111001",
765=>"1111110101010001",
766=>"0010011011111100",
767=>"0000011000101010",
768=>"1101100011001111",
769=>"1110110110111010",
770=>"0000101101010000",
771=>"0001011000100110",
772=>"1111010011101101",
773=>"1011011010001100",
774=>"1111011010111101",
775=>"0111010101110100",
776=>"0100111001101011",
777=>"1101011000010101",
778=>"1011101011101001",
779=>"1110110111011001",
780=>"0010001010101100",
781=>"0001010000111101",
782=>"1101110111111110",
783=>"1110010001011010",
784=>"0000011011111011",
785=>"0001010110001111",
786=>"0000001000110110",
787=>"1011111100001101",
788=>"1101100100110011",
789=>"0110000100010111",
790=>"0110011110001000",
791=>"1110110011010000",
792=>"1011011110100111",
793=>"1101111011100011",
794=>"0001100111001110",
795=>"0001111110010000",
796=>"1110100000001011",
797=>"1101110101001111",
798=>"0000000010000010",
799=>"0001010000000010",
800=>"0000110001101000",
801=>"1100111000000000",
802=>"1100001011011010",
803=>"0100001111011101",
804=>"0111100010001100",
805=>"0000101010101101",
806=>"1011101011101011",
807=>"1100111011010010",
808=>"0000110100001111",
809=>"0010010110011001",
810=>"1111011100100010",
811=>"1101100000100000",
812=>"1111011100000011",
813=>"0000111111001100",
814=>"0001010010011110",
815=>"1110001001100101",
816=>"1011011001110011",
817=>"0001101110101011",
818=>"0111111010001011",
819=>"0010111011100010",
820=>"1100010000000011",
821=>"1100001110011111",
822=>"1111111001110110",
823=>"0010011100110010",
824=>"0000010011111011",
825=>"1101100010111100",
826=>"1110110111111011",
827=>"0000110000001011",
828=>"0001011000001011",
829=>"1111001111000100",
830=>"1011011011010100",
831=>"1111100011110001",
832=>"0111011000001111",
833=>"0100110001000111",
834=>"1101010010110000",
835=>"1011101100001001",
836=>"1110111011001001",
837=>"0010001011010010",
838=>"0001001101011111",
839=>"1101110111010100",
840=>"1110010010111001",
841=>"0000011100010011",
842=>"0001010110101110",
843=>"0000000110100100",
844=>"1011111100100001",
845=>"1101101100110010",
846=>"0110000111101001",
847=>"0110011010001111",
848=>"1110101100110100",
849=>"1011011011111110",
850=>"1101111101011000",
851=>"0001101011101100",
852=>"0001111010101101",
853=>"1110011110000111",
854=>"1101110110011110",
855=>"0000000010011000",
856=>"0001001110010000",
857=>"0000110000100111",
858=>"1100110101010110",
859=>"1100010000100001",
860=>"0100010010111000",
861=>"0111011111010110",
862=>"0000011111111101",
863=>"1011100101101100",
864=>"1101000110111110",
865=>"0000111111110100",
866=>"0010010010011000",
867=>"1111010000001100",
868=>"1101100010111111",
869=>"1111100011101000",
870=>"0001000011001001",
871=>"0001001100001011",
872=>"1101111001011110",
873=>"1011100000001010",
874=>"0010001101110001",
875=>"0111111010100101",
876=>"0010011110110100",
877=>"1100000111010001",
878=>"1100010111100101",
879=>"0000001000010101",
880=>"0010011110100110",
881=>"0000000111100000",
882=>"1101100000101111",
883=>"1110111111001000",
884=>"0000110110000110",
885=>"0001011000011001",
886=>"1110111110110111",
887=>"1011010101111110",
888=>"0000000001001100",
889=>"0111100010100111",
890=>"0100011010011111",
891=>"1101000000001001",
892=>"1011110010010110",
893=>"1111001001100111",
894=>"0010010001001100",
895=>"0001000010010011",
896=>"1101110011010010",
897=>"1110011011011110",
898=>"0000100010110011",
899=>"0001011000100001",
900=>"1111111011000001",
901=>"1011110000110101",
902=>"1110000100100110",
903=>"0110011110010000",
904=>"0110000101011001",
905=>"1110011000001000",
906=>"1011011111100111",
907=>"1110001110001000",
908=>"0001110101010111",
909=>"0001101110110000",
910=>"1110010011010001",
911=>"1101111010111110",
912=>"0000000101011110",
913=>"0001010001101010",
914=>"0000101110001111",
915=>"1100110001110010",
916=>"1100010111101110",
917=>"0100011011110001",
918=>"0111011110011100",
919=>"0000011011000101",
920=>"1011100100000100",
921=>"1101001010010010",
922=>"0001000000011001",
923=>"0010010011000111",
924=>"1111001101011010",
925=>"1101100111000101",
926=>"1111100100100010",
927=>"0001000010101000",
928=>"0001001011101111",
929=>"1101110111111011",
930=>"1011011111111010",
931=>"0010010101000010",
932=>"0111111010010111",
933=>"0010010110111010",
934=>"1100000011101111",
935=>"1100011000111011",
936=>"0000000111111001",
937=>"0010011101010101",
938=>"0000000111001001",
939=>"1101011111001011",
940=>"1111000001111000",
941=>"0000110110001001",
942=>"0001010101111001",
943=>"1110111010001110",
944=>"1011010100100100",
945=>"0000001001010110",
946=>"0111100110110001",
947=>"0100010001100010",
948=>"1100111100000001",
949=>"1011110110001010",
950=>"1111001010101000",
951=>"0010010010100010",
952=>"0001000001101010",
953=>"1101101111101011",
954=>"1110011110011111",
955=>"0000100011101111",
956=>"0001011000010100",
957=>"1111110111000101",
958=>"1011101110011010",
959=>"1110000111100011",
960=>"0110100001100010",
961=>"0110000000001110",
962=>"1110010010110100",
963=>"1011011110110001",
964=>"1110010000001111",
965=>"0001110111000001",
966=>"0001101110001110",
967=>"1110010010111101",
968=>"1101111110011110",
969=>"0000001001000001",
970=>"0001001110100000",
971=>"0000100110110011",
972=>"1100100011111011",
973=>"1100100110110111",
974=>"0100111000010001",
975=>"0111001110100110",
976=>"1111111110110101",
977=>"1011100011110111",
978=>"1101010110100001",
979=>"0001001100110001",
980=>"0010001101110000",
981=>"1111000001001000",
982=>"1101100111001101",
983=>"1111101101011001",
984=>"0001000100001101",
985=>"0001000101110110",
986=>"1101100101101011",
987=>"1011101011111101",
988=>"0010110101100010",
989=>"0111110111000001",
990=>"0001111010110110",
991=>"1011111000010110",
992=>"1100100101100110",
993=>"0000010100001001",
994=>"0010011101111011",
995=>"1111111011011001",
996=>"1101011111111011",
997=>"1111001010001001",
998=>"0000110111111111",
999=>"0001010101111101",
1000=>"1110101100010000",
1001=>"1011010100101100",
1002=>"0000100110101101",
1003=>"0111101100111001",
1004=>"0011110110011110",
1005=>"1100101110101100",
1006=>"1011111100001001",
1007=>"1111011001011101",
1008=>"0010010101011010",
1009=>"0000110001011001",
1010=>"1101101011100111",
1011=>"1110100101001111",
1012=>"0000101000110100",
1013=>"0001011001010001",
1014=>"1111101010101110",
1015=>"1011101000110111",
1016=>"1110100100110000",
1017=>"0110110101010001",
1018=>"0101101100101101",
1019=>"1110001100110010",
1020=>"1011100001011110",
1021=>"1110010011110110",
1022=>"0001111010000101",
1023=>"0001101001001001");
  
  rom5 <= (
0=>"1110001111100110",
1=>"1101111110001010",
2=>"0000001100100010",
3=>"0001010001100111",
4=>"0000100110011011",
5=>"1100011110011111",
6=>"1100101100100100",
7=>"0100111111011000",
8=>"0111001110000000",
9=>"1111111010000011",
10=>"1011100001111001",
11=>"1101011001011101",
12=>"0001010001110000",
13=>"0010001100110100",
14=>"1110111100110111",
15=>"1101100111010110",
16=>"1111101110100000",
17=>"0001001001100100",
18=>"0001000101101010",
19=>"1101100000111111",
20=>"1011101100000111",
21=>"0010111011001010",
22=>"0111110110011100",
23=>"0001110011101111",
24=>"1011110101111110",
25=>"1100100101100110",
26=>"0000011001010011",
27=>"0010011011101110",
28=>"1111111000001000",
29=>"1101100000111000",
30=>"1111001100010010",
31=>"0000111011011001",
32=>"0001010101000010",
33=>"1110100111011000",
34=>"1011010110001101",
35=>"0000101110101101",
36=>"0111101110001001",
37=>"0011110001011100",
38=>"1100101001100110",
39=>"1011111110000000",
40=>"1111011111101001",
41=>"0010010111100000",
42=>"0000101110001110",
43=>"1101101001010101",
44=>"1110100111011100",
45=>"0000100111010100",
46=>"0001011001111001",
47=>"1111101011010000",
48=>"1011100011000100",
49=>"1110101100010010",
50=>"0110111010011111",
51=>"0101100110001100",
52=>"1101111000110001",
53=>"1011100100010010",
54=>"1110100001110111",
55=>"0010000001000001",
56=>"0001100001011000",
57=>"1110000111101010",
58=>"1110000101100110",
59=>"0000010001101000",
60=>"0001010011110011",
61=>"0000011101001000",
62=>"1100010011111111",
63=>"1100111111101111",
64=>"0101011001110100",
65=>"0110111100010001",
66=>"1111011110000011",
67=>"1011011110111000",
68=>"1101100111010100",
69=>"0001010111001111",
70=>"0010000111000110",
71=>"1110110011010101",
72=>"1101101010110010",
73=>"1111110101001110",
74=>"0001001010011100",
75=>"0000111110011110",
76=>"1101010010101001",
77=>"1011111001001111",
78=>"0011011010000001",
79=>"0111110000110100",
80=>"0001010111011111",
81=>"1011110000101001",
82=>"1100110011010101",
83=>"0000100100101110",
84=>"0010011100001110",
85=>"1111101010110001",
86=>"1101100000100001",
87=>"1111010100001100",
88=>"0000111100010100",
89=>"0001010001001100",
90=>"1110011001010000",
91=>"1011011010010011",
92=>"0001001011000110",
93=>"0111110101101000",
94=>"0011010100010111",
95=>"1100011101011110",
96=>"1100000100111000",
97=>"1111101101100011",
98=>"0010011001110000",
99=>"0000100001100110",
100=>"1101100110001111",
101=>"1110101010111000",
102=>"0000100110011010",
103=>"0001010110000011",
104=>"1111100101100101",
105=>"1011100100010110",
106=>"1110110001000110",
107=>"0110111110010111",
108=>"0101011011100111",
109=>"1101110101001011",
110=>"1011100111010001",
111=>"1110100100110100",
112=>"0010000010011011",
113=>"0001011110110001",
114=>"1110000100000110",
115=>"1110001000000101",
116=>"0000010010100111",
117=>"0001010001111010",
118=>"0000011010000101",
119=>"1100001111001010",
120=>"1101000110110000",
121=>"0101011100110000",
122=>"0110111001111101",
123=>"1111011001100110",
124=>"1011100000101000",
125=>"1101101001011110",
126=>"0001011001110001",
127=>"0010000111111011",
128=>"1110110000111101",
129=>"1101101101010000",
130=>"1111110110111010",
131=>"0001001010011011",
132=>"0000111110100110",
133=>"1101001101110010",
134=>"1011111001010110",
135=>"0011100000111100",
136=>"0111101101101100",
137=>"0001001111010111",
138=>"1011101111011111",
139=>"1100110011000101",
140=>"0000100111101111",
141=>"0010011000100001",
142=>"1111100101110111",
143=>"1101100000111010",
144=>"1111010101111011",
145=>"0001000000010101",
146=>"0001010001000101",
147=>"1110010100101001",
148=>"1011011010001100",
149=>"0001010101110100",
150=>"0111110111101011",
151=>"0011010000010011",
152=>"1100011001100110",
153=>"1100000111101111",
154=>"1111101110110000",
155=>"0010011010111001",
156=>"0000011111010101",
157=>"1101100111100110",
158=>"1110110010101110",
159=>"0000101011010011",
160=>"0001011000110110",
161=>"1111011010001000",
162=>"1011011110110000",
163=>"1111010001110100",
164=>"0111001011000100",
165=>"0101000110010001",
166=>"1101100001000010",
167=>"1011101001100000",
168=>"1110110000011101",
169=>"0010001000000000",
170=>"0001010110000100",
171=>"1101111011101110",
172=>"1110001101100000",
173=>"0000011001100101",
174=>"0001010101011110",
175=>"0000001110011000",
176=>"1100000001011100",
177=>"1101011001101110",
178=>"0101111000111001",
179=>"0110100111100111",
180=>"1110111110101001",
181=>"1011011110100001",
182=>"1101110101000010",
183=>"0001100010110100",
184=>"0010000001101101",
185=>"1110100101101100",
186=>"1101110010001110",
187=>"1111111111010010",
188=>"0001001110011010",
189=>"0000110101111001",
190=>"1100111110001001",
191=>"1100001000001010",
192=>"0011111110100100",
193=>"0111100110101100",
194=>"0000110100111111",
195=>"1011101001101110",
196=>"1101000001010001",
197=>"0000110110001100",
198=>"0010010111000001",
199=>"1111011011000000",
200=>"1101100011010001",
201=>"1111011101011010",
202=>"0000111110001000",
203=>"0001001100011100",
204=>"1110000110011010",
205=>"1011011100000111",
206=>"0001110101001100",
207=>"0111111011100101",
208=>"0011000111011011",
209=>"1100011010001001",
210=>"1100001001001000",
211=>"1111110100001100",
212=>"0010011011000011",
213=>"0000011101000001",
214=>"1101100101010001",
215=>"1110110011101000",
216=>"0000101110010111",
217=>"0001011000010101",
218=>"1111010110000100",
219=>"1011011101011000",
220=>"1111010101100111",
221=>"0111010001100100",
222=>"0100111101110100",
223=>"1101011011000000",
224=>"1011101011110010",
225=>"1110110110001101",
226=>"0010000111110010",
227=>"0001010011010100",
228=>"1101111010010111",
229=>"1110001111100011",
230=>"0000011001011101",
231=>"0001010110011100",
232=>"0000001011101101",
233=>"1100000001111111",
234=>"1101100001001001",
235=>"0101111100111101",
236=>"0110100011000111",
237=>"1110111011110100",
238=>"1011100010000000",
239=>"1101111010010010",
240=>"0001100110100000",
241=>"0001111111000001",
242=>"1110100010110010",
243=>"1101110100001011",
244=>"1111111110110110",
245=>"0001001101100111",
246=>"0000110011100100",
247=>"1100111101111010",
248=>"1100001011101001",
249=>"0100000100001010",
250=>"0111100100101100",
251=>"0000101101000101",
252=>"1011101000000000",
253=>"1101000001001100",
254=>"0000111010001001",
255=>"0010010100011001",
256=>"1111010110000111",
257=>"1101100010000001",
258=>"1111011111110001",
259=>"0001000001110011",
260=>"0001001101111001",
261=>"1110000001011100",
262=>"1011011100111111",
263=>"0001111110100011",
264=>"0111111010010100",
265=>"0010101100110110",
266=>"1100001100001101",
267=>"1100010011010101",
268=>"0000000001011010",
269=>"0010011110111101",
270=>"0000001101000001",
271=>"1101100011110000",
272=>"1110111100111000",
273=>"0000110011101011",
274=>"0001011001001100",
275=>"1111000110000000",
276=>"1011010111001110",
277=>"1111110010100110",
278=>"0111011101000001",
279=>"0100100111100111",
280=>"1101000111110110",
281=>"1011110001011001",
282=>"1111000100110000",
283=>"0010001110001010",
284=>"0001001000010101",
285=>"1101110101111010",
286=>"1110010111111101",
287=>"0000100000001010",
288=>"0001011000010111",
289=>"0000000000101000",
290=>"1011110101101100",
291=>"1101111000001010",
292=>"0110010001001001",
293=>"0110001111100111",
294=>"1110100011001010",
295=>"1011011110100101",
296=>"1110000111101011",
297=>"0001110001001011",
298=>"0001110011001110",
299=>"1110010111101001",
300=>"1101111000110000",
301=>"0000000101010100",
302=>"0001010000011010",
303=>"0000110000100100",
304=>"1100101100111001",
305=>"1100011101010100",
306=>"0100100011111111",
307=>"0111011000010001",
308=>"0000010101011011",
309=>"1011100101010000",
310=>"1101001101000101",
311=>"0001000101011001",
312=>"0010010001001000",
313=>"1111001011100000",
314=>"1101100100010101",
315=>"1111100001011111",
316=>"0001000000100101",
317=>"0001001110010110",
318=>"1101111110101001",
319=>"1011100001101001",
320=>"0010000111011010",
321=>"0111110111000111",
322=>"0010100101101001",
323=>"1100001000010001",
324=>"1100010100101001",
325=>"0000000001010010",
326=>"0010011101001100",
327=>"0000001101100100",
328=>"1101100011000101",
329=>"1110111101101101",
330=>"0000110100010011",
331=>"0001010110101110",
332=>"1111000000111101",
333=>"1011010111011111",
334=>"1111111100100101",
335=>"0111100000111011",
336=>"0100011111000000",
337=>"1101000011101011",
338=>"1011110011010101",
339=>"1111000011110100",
340=>"0010010000010011",
341=>"0001000111010011",
342=>"1101110010100110",
343=>"1110011010100100",
344=>"0000100001011100",
345=>"0001011000000001",
346=>"1111111100110111",
347=>"1011110011010011",
348=>"1101111110010010",
349=>"0110010111010001",
350=>"0110001010101001",
351=>"1110011110001001",
352=>"1011100001001100",
353=>"1110001011111111",
354=>"0001110011000101",
355=>"0001110010011011",
356=>"1110010111101011",
357=>"1101111011011010",
358=>"0000000110001101",
359=>"0001001101011100",
360=>"0000101010111000",
361=>"1100101010101110",
362=>"1100011110001111",
363=>"0100101010111001",
364=>"0111010100111000",
365=>"0000001110110111",
366=>"1011100101000101",
367=>"1101010011001010",
368=>"0001001000100011",
369=>"0010001111101010",
370=>"1111000111011010",
371=>"1101100101001110",
372=>"1111101010001101",
373=>"0001000010100011",
374=>"0001001000011011",
375=>"1101110000001000",
376=>"1011101000010101",
377=>"0010100011011011",
378=>"0111110111101000",
379=>"0010001001000010",
380=>"1011111111100101",
381=>"1100100000110001",
382=>"0000001101110110",
383=>"0010011110001011",
384=>"0000000001110000",
385=>"1101100000010000",
386=>"1111000110001010",
387=>"0000110110010011",
388=>"0001010110101100",
389=>"1110110011111010",
390=>"1011010111111000",
391=>"0000010111100111",
392=>"0111101000111100",
393=>"0100000011110001",
394=>"1100110101111101",
395=>"1011111000110100",
396=>"1111010010101100",
397=>"0010010011101111",
398=>"0000110111001000",
399=>"1101101110001001",
400=>"1110100001000111",
401=>"0000100110110010",
402=>"0001011000110111",
403=>"1111110001010010",
404=>"1011101100001010",
405=>"1110011000100010",
406=>"0110100111100011",
407=>"0101110100011010",
408=>"1110001011110111",
409=>"1011100010101110",
410=>"1110010110010100",
411=>"0001111011001001",
412=>"0001101000001000",
413=>"1110001110011110",
414=>"1110000010100011",
415=>"0000001100010101",
416=>"0001010001001000",
417=>"0000100110000101",
418=>"1100011011110110",
419=>"1100110110001001",
420=>"0101000001101001",
421=>"0111010001110111",
422=>"0000001000011111",
423=>"1011100010000001",
424=>"1101010100011100",
425=>"0001001011011110",
426=>"0010010000011011",
427=>"1111000001101000",
428=>"1101101001001010",
429=>"1111101011000010",
430=>"0001001000010100",
431=>"0001001000000010",
432=>"1101101000101100",
433=>"1011101010001111",
434=>"0010101100111001",
435=>"0111110111011111",
436=>"0010000010001010",
437=>"1011111100100000",
438=>"1100100100000011",
439=>"0000010011001000",
440=>"0010011100010100",
441=>"1111111110001100",
442=>"1101100001010110",
443=>"1111001000000011",
444=>"0000111001111010",
445=>"0001010101110001",
446=>"1110101111000111",
447=>"1011010101110101",
448=>"0000011111111010",
449=>"0111101010001100",
450=>"0011111111000001",
451=>"1100110000100111",
452=>"1011111010100101",
453=>"1111011000110001",
454=>"0010010110000110",
455=>"0000110011111110",
456=>"1101101011110000",
457=>"1110100011010101",
458=>"0000100101010010",
459=>"0001011001100101",
460=>"1111110001100001",
461=>"1011101000100010",
462=>"1110100001010111",
463=>"0110101111011111",
464=>"0101101111011101",
465=>"1110000101010000",
466=>"1011100110000010",
467=>"1110011100001001",
468=>"0001111101010101",
469=>"0001100110001010",
470=>"1110001011111000",
471=>"1110000010001101",
472=>"0000001110111110",
473=>"0001010010110011",
474=>"0000100001111000",
475=>"1100011010001000",
476=>"1100110110001011",
477=>"0101001101000000",
478=>"0111000100001001",
479=>"1111101100110010",
480=>"1011100010111110",
481=>"1101100001100111",
482=>"0001010010001011",
483=>"0010001001111111",
484=>"1110111001000110",
485=>"1101101000100100",
486=>"1111110001111101",
487=>"0001001000111101",
488=>"0001000001100011",
489=>"1101011001111011",
490=>"1011110100000011",
491=>"0011001010110100",
492=>"0111110100000010",
493=>"0001100100101101",
494=>"1011110111100111",
495=>"1100101101101110",
496=>"0000011111011011",
497=>"0010011010011110",
498=>"1111101111110110",
499=>"1101100000100100",
500=>"1111010000001111",
501=>"0000111010101000",
502=>"0001010010101000",
503=>"1110100000010110",
504=>"1011011010110100",
505=>"0000111110011100",
506=>"0111110001101001",
507=>"0011011111011100",
508=>"1100100100010010",
509=>"1100000000110011",
510=>"1111100111000000",
511=>"0010011000100001",
512=>"0000100111110101",
513=>"1101100111101110",
514=>"1110101011011111",
515=>"0000101010010101",
516=>"0001011000110011",
517=>"1111100010001001",
518=>"1011100011000110",
519=>"1110111011101100",
520=>"0111000010001100",
521=>"0101011001101011",
522=>"1101101111101010",
523=>"1011100111101010",
524=>"1110101000011000",
525=>"0010000111001110",
526=>"0001011010100111",
527=>"1110000010001101",
528=>"1110000101110111",
529=>"0000001111100000",
530=>"0001010001000101",
531=>"0000011111100011",
532=>"1100011000010001",
533=>"1100111011111100",
534=>"0101010000111101",
535=>"0111000001010001",
536=>"1111100110010110",
537=>"1011100000110001",
538=>"1101100011110001",
539=>"0001010100010111",
540=>"0010001011010110",
541=>"1110110110001111",
542=>"1101101011011011",
543=>"1111110011001101",
544=>"0001001001100011",
545=>"0001000000111010",
546=>"1101010110110010",
547=>"1011110110001000",
548=>"0011010001011000",
549=>"0111110001011010",
550=>"0001011100010100",
551=>"1011110100010011",
552=>"1100110000010010",
553=>"0000100001000000",
554=>"0010011010000000",
555=>"1111101011101111",
556=>"1101100000110101",
557=>"1111010001110000",
558=>"0000111110111011",
559=>"0001010010010010",
560=>"1110011100011000",
561=>"1011011000110101",
562=>"0001000110001110",
563=>"0111101111101010",
564=>"0011011110000011",
565=>"1100100010111110",
566=>"1100000011101000",
567=>"1111101000001000",
568=>"0010011001111001",
569=>"0000100101010101",
570=>"1101101001010100",
571=>"1110101110101100",
572=>"0000101001011011",
573=>"0001011000101101",
574=>"1111100001000010",
575=>"1011100001010000",
576=>"1111000100001001",
577=>"0111000011101001",
578=>"0101010010010100",
579=>"1101101010001111",
580=>"1011100111011111",
581=>"1110101001100010",
582=>"0010000101001101",
583=>"0001011010101010",
584=>"1110000010000111",
585=>"1110001011000010",
586=>"0000010110100000",
587=>"0001010101000010",
588=>"0000010101100110",
589=>"1100001010111110",
590=>"1101010010111011",
591=>"0101101010111001",
592=>"0110101110011001",
593=>"1111001100000011",
594=>"1011100000110111",
595=>"1101101110011101",
596=>"0001011110001010",
597=>"0010000101001010",
598=>"1110101011000011",
599=>"1101101111110001",
600=>"1111111011110111",
601=>"0001001101100100",
602=>"0000111000101000",
603=>"1101001001100100",
604=>"1100000100101010",
605=>"0011101111000111",
606=>"0111101011100110",
607=>"0001000001111011",
608=>"1011101100110100",
609=>"1100111011010100",
610=>"0000110000110000",
611=>"0010011000001101",
612=>"1111100001011110",
613=>"1101100010001011",
614=>"1111011001111110",
615=>"0000111100010111",
616=>"0001001110010001",
617=>"1110001101110011",
618=>"1011011101000000",
619=>"0001100110010110",
620=>"0111110111011001",
621=>"0011000000011111",
622=>"1100010111010010",
623=>"1100001101101001",
624=>"1111111001101110",
625=>"0010011010011001",
626=>"0000011001111010",
627=>"1101100010101100",
628=>"1110110111100111",
629=>"0000101101001001",
630=>"0001010111001011",
631=>"1111010010010010",
632=>"1011011111001000",
633=>"1111011000011011",
634=>"0111001001000011",
635=>"0101001011010011",
636=>"1101100110111011",
637=>"1011101100001111",
638=>"1110101111010111",
639=>"0010000100111010",
640=>"0001011000011110",
641=>"1101111110000001",
642=>"1110001011111011",
643=>"0000010110110111",
644=>"0001010101110110",
645=>"0000010000110111",
646=>"1100000111100101",
647=>"1101010110000010",
648=>"0101110001110000",
649=>"0110101000111101",
650=>"1111000111010011",
651=>"1011100001111000",
652=>"1101110100000101",
653=>"0001100001110101",
654=>"0001111111110010",
655=>"1110100111100001",
656=>"1101110010010111",
657=>"1111111110100011",
658=>"0001001100000101",
659=>"0000110111001110",
660=>"1101000100110000",
661=>"1100000111010010",
662=>"0011110111010111",
663=>"0111100110101110",
664=>"0000111000111010",
665=>"1011101010111101",
666=>"1100111011011001",
667=>"0000110100010111",
668=>"0010010110001100",
669=>"1111011100000101",
670=>"1101100001010011",
671=>"1111011011101110",
672=>"0001000000101100",
673=>"0001001110111110",
674=>"1110001010111101",
675=>"1011011111011000",
676=>"0001101111010111",
677=>"0111110111010011",
678=>"0010111001001110",
679=>"1100010010011011",
680=>"1100001110011100",
681=>"1111111011001111",
682=>"0010011110001111",
683=>"0000010011100110",
684=>"1101100100011101",
685=>"1110111001001011",
686=>"0000110001100001",
687=>"0001011001101001",
688=>"1111001110100010",
689=>"1011011100110001",
690=>"1111100101000101",
691=>"0111010111010001",
692=>"0100110011100000",
693=>"1101010011001101",
694=>"1011110010111011",
695=>"1110111101011100",
696=>"0010001011111110",
697=>"0001001101100100",
698=>"1101111001001111",
699=>"1110010100001010",
700=>"0000011101101001",
701=>"0001011000000011",
702=>"0000000101110110",
703=>"1011111100111110",
704=>"1101101101111000",
705=>"0110000101110110",
706=>"0110011001111011",
707=>"1110101101111110",
708=>"1011011110010011",
709=>"1110000000110000",
710=>"0001101101011010",
711=>"0001110110101110",
712=>"1110011101101001",
713=>"1101111000100010",
714=>"0000000001110111",
715=>"0001001111011100",
716=>"0000110100010010",
717=>"1100110100000111",
718=>"1100010100111001",
719=>"0100010011000011",
720=>"0111011110100101",
721=>"0000100001110001",
722=>"1011101000100100",
723=>"1101001001110010",
724=>"0000111111010100",
725=>"0010010011100100",
726=>"1111010001001100",
727=>"1101100011101111",
728=>"1111100011110001",
729=>"0001000010110000",
730=>"0001001001000111",
731=>"1101111010111100",
732=>"1011100001110000",
733=>"0010001011010010",
734=>"0111111000100101",
735=>"0010011100101010",
736=>"1100001001000110",
737=>"1100011001110101",
738=>"0000000110101000",
739=>"0010011001110110",
740=>"0000001111110100",
741=>"1101100100100101",
742=>"1110111001100111",
743=>"0000110010010000",
744=>"0001010111110000",
745=>"1111001011000001",
746=>"1011011100000010",
747=>"1111101100111000",
748=>"0111010110001010",
749=>"0100101011001111",
750=>"1101001110001110",
751=>"1011110010000100",
752=>"1110111100100110",
753=>"0010001101111100",
754=>"0001001101001000",
755=>"1101111001000001",
756=>"1110010101111101",
757=>"0000011111100111",
758=>"0001010111000101",
759=>"0000000011001110",
760=>"1011111100110100",
761=>"1101110100000111",
762=>"0110001010101101",
763=>"0110010010101111",
764=>"1110101001101000",
765=>"1011100000001011",
766=>"1110000101100101",
767=>"0001101110111001",
768=>"0001110110100110",
769=>"1110011100011100",
770=>"1101111000100100",
771=>"0000000011001100",
772=>"0001001100100010",
773=>"0000101110011100",
774=>"1100110010011110",
775=>"1100011001000100",
776=>"0100011100011001",
777=>"0111011011010101",
778=>"0000011011010011",
779=>"1011100111011000",
780=>"1101001100101111",
781=>"0001000011101110",
782=>"0010010001001000",
783=>"1111001111000101",
784=>"1101100101111111",
785=>"1111100110001000",
786=>"0001000001011010",
787=>"0001001010010111",
788=>"1101110111111011",
789=>"1011100100101000",
790=>"0010010100001101",
791=>"0111111000010001",
792=>"0010010011100101",
793=>"1100000100101110",
794=>"1100011011100001",
795=>"0000001000010100",
796=>"0010011011011111",
797=>"0000000110111011",
798=>"1101100001001010",
799=>"1111000010000000",
800=>"0000110100100110",
801=>"0001010111010111",
802=>"1110111011001111",
803=>"1011011000100000",
804=>"0000001000101101",
805=>"0111100100011111",
806=>"0100010000101111",
807=>"1100111101110100",
808=>"1011111000100001",
809=>"1111001100001000",
810=>"0010010001100001",
811=>"0000111101010000",
812=>"1101110000000101",
813=>"1110011111001100",
814=>"0000100110011100",
815=>"0001011000000010",
816=>"1111110111101100",
817=>"1011110000000010",
818=>"1110001100001000",
819=>"0110011110000110",
820=>"0101111111000001",
821=>"1110010110011010",
822=>"1011100001011110",
823=>"1110001111110001",
824=>"0001110111001110",
825=>"0001101100110100",
826=>"1110010010101001",
827=>"1101111111101101",
828=>"0000001001001100",
829=>"0001010000100001",
830=>"0000101001110011",
831=>"1100100011010100",
832=>"1100101011100100",
833=>"0100111000011101",
834=>"0111001110000001",
835=>"0000000001011100",
836=>"1011100011011101",
837=>"1101010100110110",
838=>"0001001011010010",
839=>"0010001110100110",
840=>"1111000010100111",
841=>"1101100111111010",
842=>"1111101101000101",
843=>"0001000111010100",
844=>"0001000110001010",
845=>"1101100111011100",
846=>"1011101100001101",
847=>"0010011111001001",
848=>"0111110110001001",
849=>"0010001110000111",
850=>"1100000010111110",
851=>"1100100001010001",
852=>"0000001100011010",
853=>"0010011100110000",
854=>"0000000100001111",
855=>"1101100010000010",
856=>"1111000011110001",
857=>"0000111000100001",
858=>"0001010101111110",
859=>"1110111000100110",
860=>"1011011011000110",
861=>"0000010000011011",
862=>"0111100110001100",
863=>"0100001100001111",
864=>"1100111011100000",
865=>"1011111001101111",
866=>"1111010010011011",
867=>"0010010100000010",
868=>"0000111001110101",
869=>"1101101111100100",
870=>"1110100011001101",
871=>"0000100100010110",
872=>"0001011001000101",
873=>"1111110111111011",
874=>"1011110000000110",
875=>"1110010010010111",
876=>"0110100001100011",
877=>"0101111010100010",
878=>"1110001111011110",
879=>"1011100100101110",
880=>"1110010101011111",
881=>"0001111001101110",
882=>"0001101010101001",
883=>"1110010000011001",
884=>"1101111110101111",
885=>"0000001100101010",
886=>"0001010000010011",
887=>"0000100011111101",
888=>"1100100001001111",
889=>"1100101100101100",
890=>"0100111011010010",
891=>"0111001001011000",
892=>"1111111010001000",
893=>"1011100011011001",
894=>"1101011100000100",
895=>"0001001100101101",
896=>"0010001100110110",
897=>"1111000001100000",
898=>"1101100111011110",
899=>"1111101101111000",
900=>"0001001000001010",
901=>"0001000011101101",
902=>"1101100010000011",
903=>"1011101110011110",
904=>"0010111100101011",
905=>"0111110011110110",
906=>"0001110000111110",
907=>"1011111011110101",
908=>"1100101000011100",
909=>"0000011001011110",
910=>"0010011011000000",
911=>"1111110110010101",
912=>"1101100000000111",
913=>"1111001111010011",
914=>"0000111001100100",
915=>"0001010011011111",
916=>"1110100111111100",
917=>"1011011010001101",
918=>"0000101111010100",
919=>"0111101110110000",
920=>"0011101100011111",
921=>"1100101100111011",
922=>"1011111111001101",
923=>"1111011111011010",
924=>"0010010111110001",
925=>"0000101101100000",
926=>"1101101101011011",
927=>"1110100110101001",
928=>"0000101000111110",
929=>"0001010111111100",
930=>"1111101001101010",
931=>"1011101000101010",
932=>"1110101110110110",
933=>"0110110101111100",
934=>"0101011111101011",
935=>"1101111001010011",
936=>"1011100101110110",
937=>"1110100001100101",
938=>"0010000011111101",
939=>"0001011111100111",
940=>"1110000110001101",
941=>"1110000111100101",
942=>"0000010010100110",
943=>"0001010101100001",
944=>"0000011101010011",
945=>"1100010100000000",
946=>"1101000010100101",
947=>"0101010110111001",
948=>"0110111000110100",
949=>"1111011111100100",
950=>"1011100010000111",
951=>"1101101010000101",
952=>"0001010111000110",
953=>"0010001010001010",
954=>"1110111100011010",
955=>"1101101001000110",
956=>"1111110000000100",
957=>"0001001000000000",
958=>"0001000011101100",
959=>"1101100001000100",
960=>"1011110001101101",
961=>"0011000001111001",
962=>"0111110100011100",
963=>"0001101001100111",
964=>"1011111000010000",
965=>"1100101010110011",
966=>"0000011011010011",
967=>"0010011010011000",
968=>"1111110010100001",
969=>"1101011111111100",
970=>"1111010001000001",
971=>"0000111101101010",
972=>"0001010011100000",
973=>"1110100011110110",
974=>"1011011000001000",
975=>"0000110110111110",
976=>"0111101101000001",
977=>"0011101011010001",
978=>"1100101001110110",
979=>"1100000010101100",
980=>"1111100001111001",
981=>"0010011000010000",
982=>"0000101011101110",
983=>"1101101010110100",
984=>"1110101011001010",
985=>"0000100111000000",
986=>"0001011000111100",
987=>"1111100111010010",
988=>"1011100100101100",
989=>"1110110110000110",
990=>"0110111100011101",
991=>"0101011101000100",
992=>"1101110110101111",
993=>"1011100110100010",
994=>"1110100010101000",
995=>"0010000001111110",
996=>"0001011111101011",
997=>"1110000101111100",
998=>"1110000111101011",
999=>"0000010011110001",
1000=>"0001010100001110",
1001=>"0000011011000010",
1002=>"1100010100001001",
1003=>"1101000111011000",
1004=>"0101011100110001",
1005=>"0110110101101101",
1006=>"1111011011101011",
1007=>"1011100000110110",
1008=>"1101101010101010",
1009=>"0001011010101111",
1010=>"0010000111110011",
1011=>"1110110011011011",
1012=>"1101101110100100",
1013=>"1111111011001110",
1014=>"0001001100001011",
1015=>"0000111011110001",
1016=>"1101010000111101",
1017=>"1011111110011000",
1018=>"0011100000110100",
1019=>"0111101010001000",
1020=>"0001001101111010",
1021=>"1011110000010010",
1022=>"1100110101100100",
1023=>"0000101011000100");
  
  rom6 <= (
0=>"0010011001010111",
1=>"1111100111110001",
2=>"1101100001100000",
3=>"1111010110010100",
4=>"0000111010101110",
5=>"0001001111110101",
6=>"1110010101001110",
7=>"1011011011100110",
8=>"0001010110001100",
9=>"0111110010111101",
10=>"0011001110101111",
11=>"1100011100111010",
12=>"1100001001110001",
13=>"1111110010111011",
14=>"0010011001111000",
15=>"0000011111111000",
16=>"1101100111100100",
17=>"1110110011000100",
18=>"0000101011110001",
19=>"0001010110101100",
20=>"1111011001110111",
21=>"1011100000001001",
22=>"1111001110100110",
23=>"0111001100011001",
24=>"0101000011010101",
25=>"1101011111111011",
26=>"1011101100011111",
27=>"1110110001100010",
28=>"0010000110110111",
29=>"0001010100101110",
30=>"1101111101011000",
31=>"1110001110101101",
32=>"0000010111110111",
33=>"0001010110000110",
34=>"0000001111101100",
35=>"1100001000011111",
36=>"1101001101000000",
37=>"0101100100111000",
38=>"0110110010011101",
39=>"1111010010010100",
40=>"1011100010110000",
41=>"1101101101001100",
42=>"0001011101101111",
43=>"0010000010100111",
44=>"1110101101011110",
45=>"1101101111010010",
46=>"1111111011111101",
47=>"0001001010010011",
48=>"0000111011000101",
49=>"1101001011010110",
50=>"1100000001101011",
51=>"0011100111111111",
52=>"0111101011110100",
53=>"0001000100111011",
54=>"1011110010011111",
55=>"1100111000100000",
56=>"0000101110010101",
57=>"0010010111001111",
58=>"1111100011110101",
59=>"1101100010110110",
60=>"1111010111010111",
61=>"0000111111010101",
62=>"0001010000100001",
63=>"1110010010011111",
64=>"1011011101101011",
65=>"0001011111010110",
66=>"0111110010111111",
67=>"0011000100000111",
68=>"1100011000100101",
69=>"1100001001111000",
70=>"1111110101000011",
71=>"0010011100110110",
72=>"0000011100001111",
73=>"1101100111001001",
74=>"1110110100111110",
75=>"0000101111000010",
76=>"0001010110110000",
77=>"1111010110011010",
78=>"1011011110000010",
79=>"1111010111111100",
80=>"0111001100101010",
81=>"0100111100100011",
82=>"1101011100111000",
83=>"1011101111101101",
84=>"1110110111011011",
85=>"0010001000101001",
86=>"0001010011100001",
87=>"1101111011110001",
88=>"1110010010101101",
89=>"0000011100111011",
90=>"0001010110110111",
91=>"0000001100000100",
92=>"1100000101000111",
93=>"1101100001111010",
94=>"0101111011100000",
95=>"0110011111110101",
96=>"1110111011100000",
97=>"1011100001001110",
98=>"1101111011011000",
99=>"0001100101011010",
100=>"0001111011000011",
101=>"1110100010001000",
102=>"1101110110100010",
103=>"0000000001100111",
104=>"0001001110001001",
105=>"0000110111101110",
106=>"1100111101111010",
107=>"1100001110101101",
108=>"0100000010100100",
109=>"0111100001111111",
110=>"0000101111101010",
111=>"1011101010010011",
112=>"1101000100100001",
113=>"0000111001010011",
114=>"0010010101110110",
115=>"1111010110110111",
116=>"1101100011000010",
117=>"1111011111101010",
118=>"0001000001101101",
119=>"0001001010101011",
120=>"1110000010111000",
121=>"1011011110101011",
122=>"0001111011110010",
123=>"0111110100111101",
124=>"0010101011100100",
125=>"1100001101001101",
126=>"1100010110010111",
127=>"1111111111000011",
128=>"0010011011001011",
129=>"0000010010011011",
130=>"1101100011010010",
131=>"1110111010001011",
132=>"0000110011101000",
133=>"0001010110001000",
134=>"1111001000001101",
135=>"1011011011001101",
136=>"1111110100001000",
137=>"0111011010000110",
138=>"0100100001110001",
139=>"1101001100101100",
140=>"1011110011101010",
141=>"1111000011101110",
142=>"0010001110101101",
143=>"0001010010011001",
144=>"1101111011110111",
145=>"1110010100001000",
146=>"0000011111001001",
147=>"0001010101111101",
148=>"0000001001000100",
149=>"1100000001100010",
150=>"1101101000111000",
151=>"0101111111111000",
152=>"0110011001110110",
153=>"1110110011100110",
154=>"1011100010011110",
155=>"1110000000010000",
156=>"0001101010010100",
157=>"0001111010101000",
158=>"1110100001010111",
159=>"1101110101110011",
160=>"0000000000010000",
161=>"0001001011010100",
162=>"0000110010010001",
163=>"1100111001010001",
164=>"1100010001101111",
165=>"0100001001001011",
166=>"0111011111010010",
167=>"0000101000110110",
168=>"1011101001010000",
169=>"1101000111000101",
170=>"0000111110000101",
171=>"0010010011010001",
172=>"1111010100111100",
173=>"1101100100111001",
174=>"1111100010011100",
175=>"0001000000000011",
176=>"0001001100001011",
177=>"1101111111101110",
178=>"1011100001011011",
179=>"0010000100101101",
180=>"0111110100111000",
181=>"0010100011110110",
182=>"1100001011010100",
183=>"1100010110011111",
184=>"0000000010001010",
185=>"0010011011001110",
186=>"0000001101001101",
187=>"1101100001111111",
188=>"1110111101111000",
189=>"0000110011000010",
190=>"0001010111010110",
191=>"1111000100100101",
192=>"1011011011010011",
193=>"1111111001100100",
194=>"0111011111000111",
195=>"0100011010011001",
196=>"1101000110100111",
197=>"1011110100110111",
198=>"1111000110000001",
199=>"0010001110110101",
200=>"0001000011010101",
201=>"1101110010100000",
202=>"1110011011101000",
203=>"0000100011110011",
204=>"0001011000000010",
205=>"1111111101010011",
206=>"1011110100101100",
207=>"1101111111101100",
208=>"0110010100011001",
209=>"0110001001001111",
210=>"1110100000111100",
211=>"1011100010011111",
212=>"1110001011001010",
213=>"0001110010001100",
214=>"0001110001111110",
215=>"1110010110011111",
216=>"1101111101011001",
217=>"0000000101101010",
218=>"0001010000001100",
219=>"0000101100111101",
220=>"1100101101010011",
221=>"1100100011010011",
222=>"0100100111111000",
223=>"0111010001110011",
224=>"0000001101011100",
225=>"1011101000011001",
226=>"1101010010111111",
227=>"0001000100101001",
228=>"0010010001111100",
229=>"1111000111101110",
230=>"1101100111000000",
231=>"1111101000110111",
232=>"0001000110100100",
233=>"0001000111110110",
234=>"1101110010010110",
235=>"1011101001100001",
236=>"0010100100101010",
237=>"0111110011100100",
238=>"0010001001001001",
239=>"1100000001000001",
240=>"1100100001000001",
241=>"0000001111100011",
242=>"0010011101110011",
243=>"0000000011100011",
244=>"1101100010000011",
245=>"1111001000111110",
246=>"0000111010011010",
247=>"0001010011111101",
248=>"1110110101000001",
249=>"1011010111111111",
250=>"0000000011110011",
251=>"0111011101001001",
252=>"0100010101101001",
253=>"1101000101010101",
254=>"1011111001000010",
255=>"1111001001101100",
256=>"0010010000000001",
257=>"0000111111101000",
258=>"1101110010010101",
259=>"1110011111000110",
260=>"0000100010011010",
261=>"0001011000010111",
262=>"1111111110001101",
263=>"1011110100001001",
264=>"1110000110001011",
265=>"0110011000000011",
266=>"0110000010001011",
267=>"1110011011010010",
268=>"1011101111111100",
269=>"1110010111011010",
270=>"0001110000100111",
271=>"0001101000010110",
272=>"1110100100010000",
273=>"1110010001101101",
274=>"0000001110010101",
275=>"0001000111101011",
276=>"0000101010001011",
277=>"1101010111100010",
278=>"1101011100000010",
279=>"0011110100000110",
280=>"0101101010111110",
281=>"0000010001001001",
282=>"1100111110000011",
283=>"1110010100110000",
284=>"0000111110100000",
285=>"0001101110110010",
286=>"1111101011011001",
287=>"1110101100000000",
288=>"0000000110010111",
289=>"0000111010100101",
290=>"0000111011100011",
291=>"1110111011111001",
292=>"1101111001011111",
293=>"0001101111010110",
294=>"0100011100110000",
295=>"0001010110010101",
296=>"1110010101100001",
297=>"1110101110101101",
298=>"0000011111101010",
299=>"0001011100001100",
300=>"0000011001100111",
301=>"1111011000110000",
302=>"0000000110000011",
303=>"0000110000001011",
304=>"0000111011010011",
305=>"1111111110010110",
306=>"1110111110010101",
307=>"0000100111011100",
308=>"0010101111101000",
309=>"0001100001100001",
310=>"1111101011110101",
311=>"1111011110100011",
312=>"0000011110110001",
313=>"0000111011010011",
314=>"0000110000110100",
315=>"0000000110000111",
316=>"0000011011111101",
317=>"0000100110100011",
318=>"0000110000110001",
319=>"0000100000011111",
320=>"0000010011101011",
321=>"0000011011011111",
322=>"0001001010110001",
323=>"0000101100111010",
324=>"0000111001100111",
325=>"0000000110100111",
others=>(others=>'0'));
end architecture;
